package data14_7;
localparam logic signed [13:0] dlWeights [0:1279] = {
14'b00000000100000, 
14'b00000000000001, 
14'b11111111100111, 
14'b00000000000000, 
14'b11111111110111, 
14'b00000000010001, 
14'b00000000001000, 
14'b11111111100110, 
14'b00000000000101, 
14'b00000000010101, 
14'b00000000010101, 
14'b11111111011110, 
14'b11111111001111, 
14'b11111111101010, 
14'b00000000001100, 
14'b11111111110000, 
14'b11111111110110, 
14'b11111111111100, 
14'b11111111111001, 
14'b11111111111111, 
14'b00000000001111, 
14'b11111111100001, 
14'b00000000000110, 
14'b00000000001010, 
14'b11111111111011, 
14'b00000000000000, 
14'b11111111110111, 
14'b00000000000100, 
14'b00000000001000, 
14'b00000000100000, 
14'b00000001001001, 
14'b11111111001001, 
14'b11111111100000, 
14'b11111111011010, 
14'b11111111100010, 
14'b00000000001111, 
14'b11111111111100, 
14'b00000000010100, 
14'b11111111110110, 
14'b00000000011010, 
14'b00000000010011, 
14'b11111111101110, 
14'b11111111111101, 
14'b11111111101010, 
14'b00000000000000, 
14'b11111111110011, 
14'b00000000010110, 
14'b11111111101100, 
14'b11111111110001, 
14'b00000000000001, 
14'b00000000101110, 
14'b11111111101101, 
14'b11111111011111, 
14'b11111111010101, 
14'b11111111101011, 
14'b00000000001100, 
14'b11111111111101, 
14'b00000000010000, 
14'b00000000001000, 
14'b00000000001101, 
14'b00000000011111, 
14'b11111111100110, 
14'b00000000001000, 
14'b00000000001000, 
14'b11111111101010, 
14'b00000000011101, 
14'b00000000011011, 
14'b00000000000000, 
14'b00000000010110, 
14'b11111111110101, 
14'b00000000000000, 
14'b00000000011010, 
14'b11111111100011, 
14'b11111111101100, 
14'b11111111101011, 
14'b00000000001100, 
14'b11111111111010, 
14'b00000000010110, 
14'b11111111100010, 
14'b11111111101000, 
14'b11111111110110, 
14'b11111111110010, 
14'b11111111100011, 
14'b00000000001101, 
14'b11111111101110, 
14'b00000000010001, 
14'b00000000000000, 
14'b11111111101010, 
14'b11111111111000, 
14'b11111111110001, 
14'b00000000000100, 
14'b00000000000010, 
14'b11111111110010, 
14'b00000000000011, 
14'b11111111011100, 
14'b11111111111001, 
14'b11111111100001, 
14'b00000000101000, 
14'b11111111011110, 
14'b11111111011001, 
14'b00000000000010, 
14'b00000000100110, 
14'b00000000000000, 
14'b00000000000100, 
14'b11111111101100, 
14'b11111111111100, 
14'b11111111101001, 
14'b11111111101010, 
14'b00000000001101, 
14'b11111111100111, 
14'b00000000000011, 
14'b00000000010101, 
14'b00000000000100, 
14'b00000000010000, 
14'b11111111100000, 
14'b11111111110011, 
14'b11111111011110, 
14'b00000000001110, 
14'b11111111101010, 
14'b00000000001000, 
14'b11111111101000, 
14'b11111111111000, 
14'b00000000000010, 
14'b00000000001001, 
14'b11111111100001, 
14'b11111111110111, 
14'b11111111100010, 
14'b11111111110011, 
14'b00000000000000, 
14'b00000000001010, 
14'b11111111101011, 
14'b11111111110111, 
14'b11111111110010, 
14'b00000000100011, 
14'b11111111101001, 
14'b11111111010111, 
14'b11111111101101, 
14'b00000000101000, 
14'b11111111111001, 
14'b00000000000110, 
14'b11111111111110, 
14'b11111111110101, 
14'b00000000000001, 
14'b00000000000110, 
14'b00000000011001, 
14'b11111111111010, 
14'b11111111011110, 
14'b00000000011010, 
14'b11111111111001, 
14'b00000000001000, 
14'b00000000000010, 
14'b00000000001010, 
14'b00000000010010, 
14'b11111111111110, 
14'b00000000001010, 
14'b11111111101101, 
14'b11111110011111, 
14'b00000000011001, 
14'b11111111111010, 
14'b00000000001100, 
14'b00000000010100, 
14'b11111111111000, 
14'b11111111011110, 
14'b00000000010111, 
14'b00000000011011, 
14'b11111111110010, 
14'b00000000100000, 
14'b11111111111000, 
14'b00000000000101, 
14'b11111111111101, 
14'b00000000010010, 
14'b11111111111110, 
14'b11111111111000, 
14'b11111111010100, 
14'b00000000000010, 
14'b00000000000111, 
14'b11111111110101, 
14'b11111111111100, 
14'b11111111110001, 
14'b00000000010010, 
14'b00000000011110, 
14'b11111111100010, 
14'b11111111111101, 
14'b11111111110100, 
14'b00000000011110, 
14'b11111111111110, 
14'b00000000010001, 
14'b11111111110001, 
14'b00000000011001, 
14'b00000000000000, 
14'b00000000011110, 
14'b11111111010011, 
14'b11111111101101, 
14'b11111111011110, 
14'b11111111111111, 
14'b00000000001011, 
14'b00000000000101, 
14'b00000000001101, 
14'b00000000010011, 
14'b11111111111010, 
14'b00000000011010, 
14'b11111111011110, 
14'b11111111110010, 
14'b11111111101110, 
14'b11111111111111, 
14'b00000000000001, 
14'b00000000000000, 
14'b11111111111011, 
14'b00000000000010, 
14'b11111111110011, 
14'b11111111111000, 
14'b11111111111010, 
14'b11111111111010, 
14'b11111111100101, 
14'b11111111111110, 
14'b00000000000011, 
14'b00000000011010, 
14'b11111111110100, 
14'b00000000000001, 
14'b00000000000101, 
14'b11111111101110, 
14'b11111111111001, 
14'b11111111100111, 
14'b00000000010111, 
14'b11111111100110, 
14'b00000000011110, 
14'b11111111101001, 
14'b00000000000010, 
14'b11111111110101, 
14'b11111111011101, 
14'b00000000010100, 
14'b00000000011101, 
14'b11111111100111, 
14'b00000000001000, 
14'b11111111111101, 
14'b00000000000001, 
14'b11111111110010, 
14'b00000000010100, 
14'b00000000000111, 
14'b00000000000110, 
14'b00000000000000, 
14'b11111111110010, 
14'b00000000001010, 
14'b00000000001111, 
14'b00000000001010, 
14'b11111111110101, 
14'b11111111101010, 
14'b11111111110111, 
14'b00000000001111, 
14'b11111111101101, 
14'b00000000001001, 
14'b00000000001000, 
14'b11111111110110, 
14'b11111111101111, 
14'b11111111011110, 
14'b11111111110010, 
14'b00000000000001, 
14'b00000000000000, 
14'b11111111011001, 
14'b11111111100101, 
14'b11111111100000, 
14'b00000000000101, 
14'b00000000000011, 
14'b00000000001011, 
14'b11111111010101, 
14'b00000000000010, 
14'b00000000001110, 
14'b11111111100101, 
14'b00000000000001, 
14'b11111111111100, 
14'b00000000000011, 
14'b00000000010111, 
14'b00000000000110, 
14'b00000000000011, 
14'b11111111111011, 
14'b11111111100110, 
14'b11111111100011, 
14'b00000000100001, 
14'b11111111011100, 
14'b00000000000010, 
14'b11111111111110, 
14'b00000000000001, 
14'b00000000001011, 
14'b11111111111001, 
14'b00000000000100, 
14'b11111111110010, 
14'b00000000001101, 
14'b11111111111111, 
14'b00000000010010, 
14'b00000000001011, 
14'b11111111110010, 
14'b00000000001110, 
14'b00000000001110, 
14'b00000000000000, 
14'b00000000001011, 
14'b11111111110011, 
14'b11111111011001, 
14'b11111111111101, 
14'b11111111101010, 
14'b11111111110111, 
14'b00000000000100, 
14'b00000000011001, 
14'b00000000000110, 
14'b00000000001011, 
14'b11111111110111, 
14'b00000000000101, 
14'b00000000001010, 
14'b11111111110111, 
14'b00000000001100, 
14'b00000000011001, 
14'b00000000001111, 
14'b00000000001001, 
14'b11111111111011, 
14'b00000000000110, 
14'b00000000010010, 
14'b00000000001010, 
14'b11111111100001, 
14'b00000000000010, 
14'b11111111111010, 
14'b11111111111111, 
14'b00000000010000, 
14'b11111111011101, 
14'b11111111101110, 
14'b00000000001101, 
14'b00000000011011, 
14'b00000000000010, 
14'b00000000011011, 
14'b11111111011111, 
14'b00000000000001, 
14'b00000000001111, 
14'b00000000100011, 
14'b11111111011110, 
14'b11111111110101, 
14'b11111111010111, 
14'b11111111111000, 
14'b00000000001100, 
14'b11111111101111, 
14'b00000000000101, 
14'b11111111110100, 
14'b11111111101101, 
14'b00000000001111, 
14'b11111111110101, 
14'b11111111111001, 
14'b11111111101000, 
14'b00000000000100, 
14'b11111111110111, 
14'b00000000000111, 
14'b11111111110010, 
14'b00000000010100, 
14'b11111111101110, 
14'b00000000010100, 
14'b11111111110110, 
14'b11111111010011, 
14'b00000000000110, 
14'b00000000010011, 
14'b00000000000001, 
14'b00000000000011, 
14'b00000000000100, 
14'b00000000010100, 
14'b11111111110011, 
14'b00000000000101, 
14'b11111111100000, 
14'b00000000010000, 
14'b00000000010010, 
14'b00000000000010, 
14'b11111111110111, 
14'b00000000001010, 
14'b11111111111000, 
14'b00000000001000, 
14'b00000000000100, 
14'b00000000000000, 
14'b00000000000011, 
14'b11111111101100, 
14'b00000000000110, 
14'b11111111111010, 
14'b00000000000100, 
14'b00000000011010, 
14'b00000000010001, 
14'b11111111111101, 
14'b11111111100110, 
14'b00000000001110, 
14'b11111111100010, 
14'b11111111110111, 
14'b11111111110011, 
14'b11111111111111, 
14'b00000000010101, 
14'b11111111111001, 
14'b00000000000000, 
14'b00000000011111, 
14'b11111111111010, 
14'b11111111111010, 
14'b11111111110111, 
14'b11111111111101, 
14'b00000000010000, 
14'b11111111101001, 
14'b11111111110100, 
14'b11111111110101, 
14'b11111111100111, 
14'b11111111101111, 
14'b11111111011110, 
14'b11111111110010, 
14'b11111111110011, 
14'b11111111011111, 
14'b00000000011000, 
14'b11111111100111, 
14'b00000000001000, 
14'b11111111101010, 
14'b11111111101011, 
14'b00000000001111, 
14'b00000000000000, 
14'b11111111101001, 
14'b00000000000101, 
14'b11111111100101, 
14'b00000000010100, 
14'b00000000001001, 
14'b11111111110110, 
14'b11111111101111, 
14'b11111111110000, 
14'b00000000001100, 
14'b11111111101000, 
14'b00000000000001, 
14'b00000000010100, 
14'b00000000001011, 
14'b00000000001101, 
14'b11111111101001, 
14'b00000000011001, 
14'b00000000010011, 
14'b00000000000011, 
14'b00000000011101, 
14'b00000000000011, 
14'b11111111011100, 
14'b00000000011011, 
14'b00000000001010, 
14'b00000000010110, 
14'b11111111100011, 
14'b11111111111010, 
14'b00000000000111, 
14'b11111111101001, 
14'b11111111101100, 
14'b11111111101101, 
14'b11111111110010, 
14'b00000000011101, 
14'b00000000000001, 
14'b00000000001101, 
14'b00000000000001, 
14'b00000000011000, 
14'b00000000010111, 
14'b11111111100001, 
14'b11111111101011, 
14'b00000000010001, 
14'b11111111101111, 
14'b11111111111011, 
14'b11111111111011, 
14'b00000000010000, 
14'b00000000000110, 
14'b11111111111110, 
14'b11111111101010, 
14'b00000000010011, 
14'b11111111111001, 
14'b00000000010101, 
14'b00000000000111, 
14'b00000000001010, 
14'b11111111110111, 
14'b00000000000010, 
14'b00000000010101, 
14'b11111111111011, 
14'b11111111111110, 
14'b11111111111101, 
14'b11111111101100, 
14'b00000000100000, 
14'b00000000000100, 
14'b11111111110000, 
14'b11111111111101, 
14'b00000000000111, 
14'b11111111111010, 
14'b11111111111010, 
14'b00000000000100, 
14'b00000000011001, 
14'b00000000001110, 
14'b00000000010110, 
14'b00000000000111, 
14'b11111111101101, 
14'b00000000000101, 
14'b11111111101101, 
14'b11111111110101, 
14'b11111111110000, 
14'b00000000000000, 
14'b00000000000010, 
14'b00000000001010, 
14'b00000000000110, 
14'b00000000001000, 
14'b11111111011001, 
14'b11111111101100, 
14'b11111111111100, 
14'b00000000000011, 
14'b00000000011110, 
14'b00000000011110, 
14'b11111111011110, 
14'b11111111111011, 
14'b00000000010000, 
14'b00000000011010, 
14'b11111111011110, 
14'b11111111101101, 
14'b00000000000011, 
14'b00000000010010, 
14'b11111111110100, 
14'b11111111110111, 
14'b11111111111001, 
14'b11111111111110, 
14'b00000000011010, 
14'b00000000010101, 
14'b11111111111101, 
14'b11111111110110, 
14'b00000000010010, 
14'b00000000001001, 
14'b00000000010001, 
14'b11111111111100, 
14'b11111111110000, 
14'b11111111111000, 
14'b11111111111100, 
14'b11111111100101, 
14'b00000000000101, 
14'b11111111100110, 
14'b00000000001100, 
14'b11111111111100, 
14'b11111111111100, 
14'b00000000010000, 
14'b00000000000010, 
14'b11111111111101, 
14'b00000000001010, 
14'b00000000001000, 
14'b00000000000110, 
14'b00000000000011, 
14'b00000000001100, 
14'b11111111101111, 
14'b00000000100000, 
14'b00000000001111, 
14'b11111111011101, 
14'b00000000000010, 
14'b11111111100100, 
14'b11111111100011, 
14'b11111111011010, 
14'b11111111111001, 
14'b11111111110101, 
14'b11111111110000, 
14'b00000000001011, 
14'b00000000000010, 
14'b11111111100111, 
14'b00000000000101, 
14'b11111111110000, 
14'b11111111110010, 
14'b11111111110100, 
14'b11111111110111, 
14'b11111111110011, 
14'b00000000000010, 
14'b11111111111001, 
14'b00000000010010, 
14'b11111111110000, 
14'b00000000000110, 
14'b00000000000011, 
14'b00000000001011, 
14'b00000000011011, 
14'b00000000000000, 
14'b11111111101110, 
14'b11111111110100, 
14'b00000000001110, 
14'b00000000010001, 
14'b11111111010111, 
14'b00000000001001, 
14'b00000000000010, 
14'b11111111011101, 
14'b00000000010110, 
14'b11111111110110, 
14'b00000000000000, 
14'b11111111101101, 
14'b00000000010110, 
14'b00000000001111, 
14'b11111111010011, 
14'b00000000010001, 
14'b00000000001011, 
14'b00000000001011, 
14'b00000000100101, 
14'b00000000001010, 
14'b00000000010100, 
14'b11111111101100, 
14'b00000000000100, 
14'b11111111111000, 
14'b00000000001000, 
14'b00000000011101, 
14'b00000000001110, 
14'b11111111010111, 
14'b00000000010100, 
14'b11111111110110, 
14'b00000000000101, 
14'b11111111101111, 
14'b11111111101001, 
14'b00000000000100, 
14'b00000000001111, 
14'b00000000000111, 
14'b11111111111000, 
14'b11111111011011, 
14'b00000000001001, 
14'b00000000000011, 
14'b00000000010010, 
14'b00000000000000, 
14'b00000000000100, 
14'b00000000010011, 
14'b00000000010001, 
14'b11111111110110, 
14'b00000000001101, 
14'b11111111101111, 
14'b11111111101111, 
14'b11111111110101, 
14'b00000000010110, 
14'b11111111110000, 
14'b11111111101001, 
14'b00000000000011, 
14'b00000000001101, 
14'b00000000010001, 
14'b11111111110011, 
14'b11111111011101, 
14'b11111111011100, 
14'b00000000001111, 
14'b00000000000001, 
14'b00000000010101, 
14'b00000000010001, 
14'b00000000001110, 
14'b00000000010111, 
14'b11111111110100, 
14'b11111111111110, 
14'b00000000000101, 
14'b00000000001001, 
14'b00000000010011, 
14'b00000000010101, 
14'b00000000011010, 
14'b11111111101111, 
14'b00000000000000, 
14'b00000000011010, 
14'b00000000010011, 
14'b00000000010010, 
14'b11111111111110, 
14'b11111111101011, 
14'b11111111111010, 
14'b11111111111011, 
14'b11111111101111, 
14'b11111111100000, 
14'b00000000010000, 
14'b00000000001111, 
14'b00000000010100, 
14'b00000000000000, 
14'b11111111110011, 
14'b11111111111010, 
14'b11111111110000, 
14'b00000000000011, 
14'b00000000000000, 
14'b00000000010111, 
14'b00000000001010, 
14'b11111111011100, 
14'b11111111101101, 
14'b11111111101001, 
14'b11111111111111, 
14'b11111111100011, 
14'b11111111111001, 
14'b11111111110110, 
14'b00000000000110, 
14'b00000000000001, 
14'b00000000000100, 
14'b11111111011001, 
14'b11111111111110, 
14'b00000000010001, 
14'b00000000011011, 
14'b11111111111101, 
14'b11111111100001, 
14'b00000000001111, 
14'b11111111111000, 
14'b00000000010110, 
14'b11111111111111, 
14'b11111111011011, 
14'b11111111110100, 
14'b00000000000010, 
14'b11111111100010, 
14'b11111111111101, 
14'b00000000010110, 
14'b11111111110110, 
14'b11111111111110, 
14'b00000000010101, 
14'b00000000000111, 
14'b11111111110110, 
14'b00000000010111, 
14'b11111111110111, 
14'b00000000001001, 
14'b00000000000001, 
14'b11111111100111, 
14'b00000000010100, 
14'b11111111110011, 
14'b00000000000001, 
14'b00000000000010, 
14'b11111111110100, 
14'b11111111111001, 
14'b00000000001110, 
14'b00000000000000, 
14'b00000000000101, 
14'b00000000001001, 
14'b11111111110001, 
14'b00000000000111, 
14'b11111111101010, 
14'b11111111111111, 
14'b11111111110011, 
14'b11111111110010, 
14'b11111111101100, 
14'b00000000000011, 
14'b00000000001010, 
14'b00000000000101, 
14'b11111111110110, 
14'b11111111101101, 
14'b00000000010101, 
14'b11111111110011, 
14'b00000000000000, 
14'b00000000011001, 
14'b00000000000000, 
14'b11111111100110, 
14'b00000000010001, 
14'b11111111101110, 
14'b00000000001011, 
14'b00000000000111, 
14'b00000000001000, 
14'b00000000010000, 
14'b11111111101100, 
14'b00000000000110, 
14'b11111111110011, 
14'b11111111101000, 
14'b00000000001101, 
14'b11111111100111, 
14'b00000000010110, 
14'b00000000000100, 
14'b11111111110111, 
14'b11111111100110, 
14'b11111111110100, 
14'b00000000010101, 
14'b11111111110000, 
14'b00000000000001, 
14'b11111111110101, 
14'b00000000011000, 
14'b11111111111011, 
14'b00000000000010, 
14'b00000000001100, 
14'b11111111110011, 
14'b11111111110001, 
14'b00000000000110, 
14'b00000000000011, 
14'b11111111100010, 
14'b00000000011011, 
14'b11111111111010, 
14'b00000000011001, 
14'b00000000001110, 
14'b00000000001100, 
14'b11111111101110, 
14'b11111111111010, 
14'b11111111111010, 
14'b11111111110111, 
14'b11111111111101, 
14'b00000000001110, 
14'b11111111110000, 
14'b00000000001100, 
14'b00000000000010, 
14'b00000000000100, 
14'b00000000001101, 
14'b00000000010100, 
14'b00000000001010, 
14'b11111111110001, 
14'b00000000000111, 
14'b11111111100001, 
14'b00000000001000, 
14'b11111111110110, 
14'b00000000001100, 
14'b11111111110100, 
14'b11111111110010, 
14'b00000000001010, 
14'b11111111101100, 
14'b11111111110011, 
14'b11111111101010, 
14'b00000000000011, 
14'b11111111110001, 
14'b00000000011100, 
14'b11111111111101, 
14'b11111111110001, 
14'b11111111111111, 
14'b00000000001010, 
14'b00000000001010, 
14'b00000000010101, 
14'b11111111110101, 
14'b11111111101000, 
14'b00000000000001, 
14'b11111111101111, 
14'b11111111110101, 
14'b11111111100100, 
14'b00000000001101, 
14'b00000000100001, 
14'b00000000001100, 
14'b00000000010100, 
14'b11111111111111, 
14'b11111111110001, 
14'b00000000010010, 
14'b11111111111000, 
14'b00000000010100, 
14'b11111111110110, 
14'b00000000000101, 
14'b11111111101000, 
14'b00000000100011, 
14'b00000000011110, 
14'b11111111110010, 
14'b11111111010111, 
14'b00000000000010, 
14'b11111111101100, 
14'b00000000100000, 
14'b11111111111100, 
14'b11111111110011, 
14'b00000000000011, 
14'b11111111110001, 
14'b11111111110010, 
14'b11111111110111, 
14'b11111111011001, 
14'b00000000000011, 
14'b11111111011010, 
14'b11111111110101, 
14'b00000000000011, 
14'b00000000001011, 
14'b11111111110001, 
14'b11111111111101, 
14'b00000000000101, 
14'b11111111110110, 
14'b11111111010101, 
14'b11111111110110, 
14'b00000000000110, 
14'b00000000000100, 
14'b00000000001001, 
14'b00000000001010, 
14'b11111111011101, 
14'b11111111110100, 
14'b00000000010110, 
14'b11111111100111, 
14'b11111111110111, 
14'b00000000011101, 
14'b11111111110011, 
14'b00000000000000, 
14'b11111111110011, 
14'b00000000000100, 
14'b11111111111010, 
14'b11111111110111, 
14'b00000000010111, 
14'b11111111100111, 
14'b11111111110111, 
14'b00000000010010, 
14'b00000000010111, 
14'b11111111111001, 
14'b00000000001000, 
14'b11111111111011, 
14'b11111111011101, 
14'b11111111110111, 
14'b00000000000100, 
14'b11111111110011, 
14'b11111111111111, 
14'b11111111111000, 
14'b11111111110011, 
14'b00000000010011, 
14'b11111111110011, 
14'b11111111110000, 
14'b00000000000001, 
14'b11111111111000, 
14'b00000000001010, 
14'b11111111101011, 
14'b00000000010100, 
14'b00000000001111, 
14'b00000000000001, 
14'b11111111111111, 
14'b11111111101110, 
14'b11111111101010, 
14'b11111111110001, 
14'b11111111110110, 
14'b11111111111011, 
14'b00000000000101, 
14'b00000000011110, 
14'b11111111110111, 
14'b11111111100011, 
14'b00000000011101, 
14'b11111111110001, 
14'b11111111111100, 
14'b00000000000100, 
14'b00000000001101, 
14'b11111111101111, 
14'b11111111110001, 
14'b11111111111001, 
14'b00000000001110, 
14'b11111111110011, 
14'b00000000001100, 
14'b00000000001110, 
14'b11111111101001, 
14'b00000000000000, 
14'b00000000000000, 
14'b11111111111001, 
14'b11111111110110, 
14'b00000000000010, 
14'b11111111111001, 
14'b00000000000111, 
14'b00000000000110, 
14'b11111111101010, 
14'b11111111110001, 
14'b00000000000011, 
14'b00000000001111, 
14'b11111111100100, 
14'b11111111011100, 
14'b11111111110011, 
14'b11111111111010, 
14'b11111111111011, 
14'b11111111111101, 
14'b11111111101101, 
14'b00000000001010, 
14'b00000000001011, 
14'b11111111110011, 
14'b00000000001101, 
14'b11111111111110, 
14'b11111111110111, 
14'b00000000010110, 
14'b11111111110000, 
14'b11111111111011, 
14'b11111111110000, 
14'b00000000000110, 
14'b00000000010010, 
14'b11111111111111, 
14'b00000000001011, 
14'b11111111011011, 
14'b00000000000011, 
14'b11111111110010, 
14'b11111111110101, 
14'b00000000010011, 
14'b11111111101000, 
14'b00000000001010, 
14'b11111111110101, 
14'b00000000000000, 
14'b00000000000000, 
14'b11111111100110, 
14'b11111111111110, 
14'b00000000000011, 
14'b11111111101101, 
14'b00000000000100, 
14'b00000000010100, 
14'b11111111110010, 
14'b00000000001111, 
14'b11111111111000, 
14'b00000000011011, 
14'b11111111010111, 
14'b11111111010110, 
14'b00000000001100, 
14'b11111111110100, 
14'b00000000000101, 
14'b11111111101110, 
14'b11111111111010, 
14'b00000000001110, 
14'b00000000000100, 
14'b11111111111111, 
14'b00000000000100, 
14'b11111111110010, 
14'b00000000010001, 
14'b11111111111111, 
14'b11111111110011, 
14'b00000000001010, 
14'b11111111111100, 
14'b00000000000001, 
14'b00000000001111, 
14'b11111111100100, 
14'b11111111110000, 
14'b11111111010111, 
14'b00000000001000, 
14'b11111111100100, 
14'b00000000001100, 
14'b00000000001001, 
14'b11111111111111, 
14'b11111111101111, 
14'b11111111110010, 
14'b00000000001110, 
14'b11111111111101, 
14'b11111111011111, 
14'b00000000011001, 
14'b11111111011100, 
14'b11111111101100, 
14'b11111111111100, 
14'b00000000000000, 
14'b11111111101001, 
14'b11111111110101, 
14'b11111111111111, 
14'b11111111111101, 
14'b11111111111010, 
14'b11111111111110, 
14'b11111111110001, 
14'b00000000011100, 
14'b11111111111000, 
14'b00000000000011, 
14'b00000000000011, 
14'b11111111111011, 
14'b00000000000101, 
14'b00000000000010, 
14'b11111111111001, 
14'b11111111111010, 
14'b00000000000110, 
14'b00000000000011, 
14'b00000000000101, 
14'b00000000001010, 
14'b11111111101101, 
14'b00000000011111, 
14'b11111111110100, 
14'b00000000000100, 
14'b11111111110101, 
14'b00000000001010, 
14'b11111111101001, 
14'b11111111101110, 
14'b11111111100011, 
14'b11111111111010, 
14'b11111111010110, 
14'b11111111111110, 
14'b11111111110001, 
14'b11111111101001, 
14'b11111111101111, 
14'b11111111110111, 
14'b11111111110001, 
14'b00000000010101, 
14'b11111111010111, 
14'b00000000100001, 
14'b11111111111010, 
14'b11111111101111, 
14'b11111111111010, 
14'b11111111100111, 
14'b00000000000100, 
14'b00000000001011, 
14'b11111111101010, 
14'b00000000000101, 
14'b11111111100010, 
14'b00000000010000, 
14'b11111111100111, 
14'b00000000000101, 
14'b11111111110100, 
14'b11111111111000, 
14'b00000000010110, 
14'b00000000010010, 
14'b11111111110011, 
14'b00000000010001, 
14'b00000000000111, 
14'b00000000000100, 
14'b00000000011011, 
14'b00000000001111, 
14'b11111111110010, 
14'b11111111110000, 
14'b00000000010111, 
14'b00000000010101, 
14'b00000000000001, 
14'b00000000001100, 
14'b00000000000101, 
14'b00000000000101, 
14'b11111111111011, 
14'b00000000010011, 
14'b11111111111100, 
14'b00000000000000, 
14'b00000000000111, 
14'b00000000100110, 
14'b11111111101010, 
14'b11111111110111, 
14'b00000000000000, 
14'b00000000010000, 
14'b00000000010011, 
14'b11111111101100, 
14'b11111111101011, 
14'b00000000000010, 
14'b00000000000111, 
14'b00000000000010, 
14'b00000000000100, 
14'b00000000001001, 
14'b00000000000111, 
14'b00000000010000, 
14'b11111111111111, 
14'b00000000000010, 
14'b00000000010010, 
14'b11111111111110, 
14'b11111111111010, 
14'b00000000000100, 
14'b11111111100110, 
14'b00000000000011, 
14'b00000000001011, 
14'b11111111101011, 
14'b00000000011111, 
14'b11111111111110, 
14'b00000000000111, 
14'b11111111111110, 
14'b11111111111011, 
14'b11111111111010, 
14'b00000000001110, 
14'b00000000011111, 
14'b00000000000000, 
14'b00000000001100, 
14'b00000000100000, 
14'b11111111100111, 
14'b00000000001111, 
14'b00000000010000, 
14'b11111111101111, 
14'b00000000000011, 
14'b00000000010011, 
14'b00000000000001, 
14'b00000000001110, 
14'b11111111111101, 
14'b00000000011011, 
14'b00000000001011, 
14'b11111111110100, 
14'b11111111100001, 
14'b11111111101101, 
14'b00000000000110, 
14'b00000000000001, 
14'b11111111111100, 
14'b00000000001000, 
14'b00000000001011, 
14'b00000000001010, 
14'b11111111100011, 
14'b00000000000101, 
14'b00000000001101, 
14'b11111111100110, 
14'b11111111110010, 
14'b11111111111011, 
14'b00000000011001, 
14'b00000000011010, 
14'b11111111111111, 
14'b00000000001110, 
14'b11111111100110, 
14'b11111111110110, 
14'b11111111110111, 
14'b11111111111100, 
14'b00000000000010, 
14'b11111111011110, 
14'b00000000001110, 
14'b11111111111001, 
14'b11111111111001, 
14'b11111111101010, 
14'b00000000000011, 
14'b11111111111110, 
14'b00000000100101, 
14'b11111111100010, 
14'b00000000001000, 
14'b00000000000000, 
14'b11111111110000, 
14'b11111111110110, 
14'b00000000000101, 
14'b11111111101010, 
14'b11111111110011, 
14'b11111111100011, 
14'b11111111111000, 
14'b00000000001101, 
14'b00000000011001, 
14'b11111111101111, 
14'b11111111111001, 
14'b00000000000100, 
14'b00000000010100, 
14'b11111111110111, 
14'b11111111111111, 
14'b11111111111101, 
14'b00000000010110, 
14'b11111111011101, 
14'b00000000010101, 
14'b11111111110010, 
14'b11111111011111, 
14'b11111111101111, 
14'b00000000100001, 
14'b11111111100101, 
14'b11111111111000, 
14'b11111111100000, 
14'b00000000001100, 
14'b00000000011100, 
14'b00000000011101, 
14'b11111111101111, 
14'b00000000000001, 
14'b11111111011110, 
14'b00000000001101, 
14'b11111111110000, 
14'b00000000010010, 
14'b00000000000000, 
14'b00000000001010, 
14'b11111111110000, 
14'b11111111110011, 
14'b11111111101110, 
14'b00000000000110, 
14'b00000000001000, 
14'b00000000011011, 
14'b00000000000100, 
14'b11111111110000, 
14'b11111111111000, 
14'b11111111100100, 
14'b00000000010101, 
14'b00000000001110, 
14'b11111111101000, 
14'b11111111111001, 
14'b11111111011110, 
14'b00000000010101, 
14'b11111111100110, 
14'b00000000011010, 
14'b11111111101111, 
14'b00000000000110, 
14'b00000000000011, 
14'b00000000010100, 
14'b11111111101101, 
14'b11111111101011, 
14'b00000000010110, 
14'b11111111110011, 
14'b00000000000010, 
14'b11111111101010, 
14'b00000000000001, 
14'b11111111110100, 
14'b00000000001110, 
14'b11111111110110, 
14'b11111111110011, 
14'b11111111110100, 
14'b00000000001100, 
14'b11111111110110, 
14'b11111111111010, 
14'b00000000001010, 
14'b00000000010011, 
14'b11111111100001, 
14'b00000000000010, 
14'b00000000000011, 
14'b11111111011111, 
14'b11111111111011, 
14'b00000000011000, 
14'b00000000001110, 
14'b11111111100011, 
14'b00000000001111, 
14'b11111111001000, 
14'b11111111100101, 
14'b11111111101001, 
14'b00000000000010, 
14'b11111111011101, 
14'b11111111110111, 
14'b00000000000010, 
14'b11111111110100, 
14'b00000000011111, 
14'b00000000000100, 
14'b00000000000001, 
14'b00000000000000, 
14'b00000000100101, 
14'b11111111101001, 
14'b11111111101011, 
14'b00000000000101, 
14'b00000000010101, 
14'b00000000010000, 
14'b00000000010000, 
14'b11111111110001, 
14'b11111111101011, 
14'b00000000000011, 
14'b11111111101110, 
14'b00000000000101, 
14'b00000000000111, 
14'b00000000000010, 
14'b11111111100010, 
14'b11111111100010, 
14'b11111111111100, 
14'b11111111111000, 
14'b11111111111011, 
14'b11111111100000, 
14'b00000000000101, 
14'b11111111110101, 
14'b11111111011010, 
14'b11111111101111, 
14'b00000000010101, 
14'b11111111100111, 
14'b00000000010010, 
14'b00000000100000, 
14'b00000000011111, 
14'b11111111111111, 
14'b11111111101010, 
14'b00000000001101, 
14'b11111111101011, 
14'b11111111110111, 
14'b00000000001100, 
14'b11111111111100, 
14'b11111111111011, 
14'b11111111111011, 
14'b00000000010000

};
localparam logic signed [13:0] dlBiases [9:0] = {
14'b00000000010101, 
14'b11111111111111, 
14'b11111111111111, 
14'b11111111111000, 
14'b11111111111000, 
14'b11111111111101, 
14'b11111111111101, 
14'b00000000001001, 
14'b11111111101000, 
14'b11111111111101

};
localparam logic signed [13:0] convWeights [0:17] = {
14'b00000000001110, 
14'b00000000111101, 
14'b11111111100001, 
14'b00000000001011, 
14'b00000000000001, 
14'b00000001000001, 
14'b00000000110011, 
14'b00000000011001, 
14'b11111111100010, 
14'b00000000101100, 
14'b11111111110100, 
14'b00000000011010, 
14'b00000000111111, 
14'b00000000010100, 
14'b00000000110001, 
14'b11111111111110, 
14'b00000000010111, 
14'b00000000001110 

};
localparam logic signed [13:0] convBiases [1:0] = {
14'b00000000000000, 
14'b00000000000000

};
endpackage