package data10_5;
localparam logic signed [9:0] dlWeights [0:1279] = {
10'b0000001000, 
10'b0000000000, 
10'b1111111001, 
10'b0000000000, 
10'b1111111101, 
10'b0000000100, 
10'b0000000010, 
10'b1111111001, 
10'b0000000001, 
10'b0000000101, 
10'b0000000101, 
10'b1111110111, 
10'b1111110011, 
10'b1111111010, 
10'b0000000011, 
10'b1111111100, 
10'b1111111101, 
10'b1111111111, 
10'b1111111110, 
10'b1111111111, 
10'b0000000011, 
10'b1111111000, 
10'b0000000001, 
10'b0000000010, 
10'b1111111110, 
10'b0000000000, 
10'b1111111101, 
10'b0000000001, 
10'b0000000010, 
10'b0000001000, 
10'b0000010010, 
10'b1111110010, 
10'b1111111000, 
10'b1111110110, 
10'b1111111000, 
10'b0000000011, 
10'b1111111111, 
10'b0000000101, 
10'b1111111101, 
10'b0000000110, 
10'b0000000100, 
10'b1111111011, 
10'b1111111111, 
10'b1111111010, 
10'b0000000000, 
10'b1111111100, 
10'b0000000101, 
10'b1111111011, 
10'b1111111100, 
10'b0000000000, 
10'b0000001011, 
10'b1111111011, 
10'b1111110111, 
10'b1111110101, 
10'b1111111010, 
10'b0000000011, 
10'b1111111111, 
10'b0000000100, 
10'b0000000010, 
10'b0000000011, 
10'b0000000111, 
10'b1111111001, 
10'b0000000010, 
10'b0000000010, 
10'b1111111010, 
10'b0000000111, 
10'b0000000110, 
10'b0000000000, 
10'b0000000101, 
10'b1111111101, 
10'b0000000000, 
10'b0000000110, 
10'b1111111000, 
10'b1111111011, 
10'b1111111010, 
10'b0000000011, 
10'b1111111110, 
10'b0000000101, 
10'b1111111000, 
10'b1111111010, 
10'b1111111101, 
10'b1111111100, 
10'b1111111000, 
10'b0000000011, 
10'b1111111011, 
10'b0000000100, 
10'b0000000000, 
10'b1111111010, 
10'b1111111110, 
10'b1111111100, 
10'b0000000001, 
10'b0000000000, 
10'b1111111100, 
10'b0000000000, 
10'b1111110111, 
10'b1111111110, 
10'b1111111000, 
10'b0000001010, 
10'b1111110111, 
10'b1111110110, 
10'b0000000000, 
10'b0000001001, 
10'b0000000000, 
10'b0000000001, 
10'b1111111011, 
10'b1111111111, 
10'b1111111010, 
10'b1111111010, 
10'b0000000011, 
10'b1111111001, 
10'b0000000000, 
10'b0000000101, 
10'b0000000001, 
10'b0000000100, 
10'b1111111000, 
10'b1111111100, 
10'b1111110111, 
10'b0000000011, 
10'b1111111010, 
10'b0000000010, 
10'b1111111010, 
10'b1111111110, 
10'b0000000000, 
10'b0000000010, 
10'b1111111000, 
10'b1111111101, 
10'b1111111000, 
10'b1111111100, 
10'b0000000000, 
10'b0000000010, 
10'b1111111010, 
10'b1111111101, 
10'b1111111100, 
10'b0000001000, 
10'b1111111010, 
10'b1111110101, 
10'b1111111011, 
10'b0000001010, 
10'b1111111110, 
10'b0000000001, 
10'b1111111111, 
10'b1111111101, 
10'b0000000000, 
10'b0000000001, 
10'b0000000110, 
10'b1111111110, 
10'b1111110111, 
10'b0000000110, 
10'b1111111110, 
10'b0000000010, 
10'b0000000000, 
10'b0000000010, 
10'b0000000100, 
10'b1111111111, 
10'b0000000010, 
10'b1111111011, 
10'b1111100111, 
10'b0000000110, 
10'b1111111110, 
10'b0000000011, 
10'b0000000101, 
10'b1111111110, 
10'b1111110111, 
10'b0000000101, 
10'b0000000110, 
10'b1111111100, 
10'b0000001000, 
10'b1111111110, 
10'b0000000001, 
10'b1111111111, 
10'b0000000100, 
10'b1111111111, 
10'b1111111110, 
10'b1111110101, 
10'b0000000000, 
10'b0000000001, 
10'b1111111101, 
10'b1111111111, 
10'b1111111100, 
10'b0000000100, 
10'b0000000111, 
10'b1111111000, 
10'b1111111111, 
10'b1111111101, 
10'b0000000111, 
10'b1111111111, 
10'b0000000100, 
10'b1111111100, 
10'b0000000110, 
10'b0000000000, 
10'b0000000111, 
10'b1111110100, 
10'b1111111011, 
10'b1111110111, 
10'b1111111111, 
10'b0000000010, 
10'b0000000001, 
10'b0000000011, 
10'b0000000100, 
10'b1111111110, 
10'b0000000110, 
10'b1111110111, 
10'b1111111100, 
10'b1111111011, 
10'b1111111111, 
10'b0000000000, 
10'b0000000000, 
10'b1111111110, 
10'b0000000000, 
10'b1111111100, 
10'b1111111110, 
10'b1111111110, 
10'b1111111110, 
10'b1111111001, 
10'b1111111111, 
10'b0000000000, 
10'b0000000110, 
10'b1111111101, 
10'b0000000000, 
10'b0000000001, 
10'b1111111011, 
10'b1111111110, 
10'b1111111001, 
10'b0000000101, 
10'b1111111001, 
10'b0000000111, 
10'b1111111010, 
10'b0000000000, 
10'b1111111101, 
10'b1111110111, 
10'b0000000101, 
10'b0000000111, 
10'b1111111001, 
10'b0000000010, 
10'b1111111111, 
10'b0000000000, 
10'b1111111100, 
10'b0000000101, 
10'b0000000001, 
10'b0000000001, 
10'b0000000000, 
10'b1111111100, 
10'b0000000010, 
10'b0000000011, 
10'b0000000010, 
10'b1111111101, 
10'b1111111010, 
10'b1111111101, 
10'b0000000011, 
10'b1111111011, 
10'b0000000010, 
10'b0000000010, 
10'b1111111101, 
10'b1111111011, 
10'b1111110111, 
10'b1111111100, 
10'b0000000000, 
10'b0000000000, 
10'b1111110110, 
10'b1111111001, 
10'b1111111000, 
10'b0000000001, 
10'b0000000000, 
10'b0000000010, 
10'b1111110101, 
10'b0000000000, 
10'b0000000011, 
10'b1111111001, 
10'b0000000000, 
10'b1111111111, 
10'b0000000000, 
10'b0000000101, 
10'b0000000001, 
10'b0000000000, 
10'b1111111110, 
10'b1111111001, 
10'b1111111000, 
10'b0000001000, 
10'b1111110111, 
10'b0000000000, 
10'b1111111111, 
10'b0000000000, 
10'b0000000010, 
10'b1111111110, 
10'b0000000001, 
10'b1111111100, 
10'b0000000011, 
10'b1111111111, 
10'b0000000100, 
10'b0000000010, 
10'b1111111100, 
10'b0000000011, 
10'b0000000011, 
10'b0000000000, 
10'b0000000010, 
10'b1111111100, 
10'b1111110110, 
10'b1111111111, 
10'b1111111010, 
10'b1111111101, 
10'b0000000001, 
10'b0000000110, 
10'b0000000001, 
10'b0000000010, 
10'b1111111101, 
10'b0000000001, 
10'b0000000010, 
10'b1111111101, 
10'b0000000011, 
10'b0000000110, 
10'b0000000011, 
10'b0000000010, 
10'b1111111110, 
10'b0000000001, 
10'b0000000100, 
10'b0000000010, 
10'b1111111000, 
10'b0000000000, 
10'b1111111110, 
10'b1111111111, 
10'b0000000100, 
10'b1111110111, 
10'b1111111011, 
10'b0000000011, 
10'b0000000110, 
10'b0000000000, 
10'b0000000110, 
10'b1111110111, 
10'b0000000000, 
10'b0000000011, 
10'b0000001000, 
10'b1111110111, 
10'b1111111101, 
10'b1111110101, 
10'b1111111110, 
10'b0000000011, 
10'b1111111011, 
10'b0000000001, 
10'b1111111101, 
10'b1111111011, 
10'b0000000011, 
10'b1111111101, 
10'b1111111110, 
10'b1111111010, 
10'b0000000001, 
10'b1111111101, 
10'b0000000001, 
10'b1111111100, 
10'b0000000101, 
10'b1111111011, 
10'b0000000101, 
10'b1111111101, 
10'b1111110100, 
10'b0000000001, 
10'b0000000100, 
10'b0000000000, 
10'b0000000000, 
10'b0000000001, 
10'b0000000101, 
10'b1111111100, 
10'b0000000001, 
10'b1111111000, 
10'b0000000100, 
10'b0000000100, 
10'b0000000000, 
10'b1111111101, 
10'b0000000010, 
10'b1111111110, 
10'b0000000010, 
10'b0000000001, 
10'b0000000000, 
10'b0000000000, 
10'b1111111011, 
10'b0000000001, 
10'b1111111110, 
10'b0000000001, 
10'b0000000110, 
10'b0000000100, 
10'b1111111111, 
10'b1111111001, 
10'b0000000011, 
10'b1111111000, 
10'b1111111101, 
10'b1111111100, 
10'b1111111111, 
10'b0000000101, 
10'b1111111110, 
10'b0000000000, 
10'b0000000111, 
10'b1111111110, 
10'b1111111110, 
10'b1111111101, 
10'b1111111111, 
10'b0000000100, 
10'b1111111010, 
10'b1111111101, 
10'b1111111101, 
10'b1111111001, 
10'b1111111011, 
10'b1111110111, 
10'b1111111100, 
10'b1111111100, 
10'b1111110111, 
10'b0000000110, 
10'b1111111001, 
10'b0000000010, 
10'b1111111010, 
10'b1111111010, 
10'b0000000011, 
10'b0000000000, 
10'b1111111010, 
10'b0000000001, 
10'b1111111001, 
10'b0000000101, 
10'b0000000010, 
10'b1111111101, 
10'b1111111011, 
10'b1111111100, 
10'b0000000011, 
10'b1111111010, 
10'b0000000000, 
10'b0000000101, 
10'b0000000010, 
10'b0000000011, 
10'b1111111010, 
10'b0000000110, 
10'b0000000100, 
10'b0000000000, 
10'b0000000111, 
10'b0000000000, 
10'b1111110111, 
10'b0000000110, 
10'b0000000010, 
10'b0000000101, 
10'b1111111000, 
10'b1111111110, 
10'b0000000001, 
10'b1111111010, 
10'b1111111011, 
10'b1111111011, 
10'b1111111100, 
10'b0000000111, 
10'b0000000000, 
10'b0000000011, 
10'b0000000000, 
10'b0000000110, 
10'b0000000101, 
10'b1111111000, 
10'b1111111010, 
10'b0000000100, 
10'b1111111011, 
10'b1111111110, 
10'b1111111110, 
10'b0000000100, 
10'b0000000001, 
10'b1111111111, 
10'b1111111010, 
10'b0000000100, 
10'b1111111110, 
10'b0000000101, 
10'b0000000001, 
10'b0000000010, 
10'b1111111101, 
10'b0000000000, 
10'b0000000101, 
10'b1111111110, 
10'b1111111111, 
10'b1111111111, 
10'b1111111011, 
10'b0000001000, 
10'b0000000001, 
10'b1111111100, 
10'b1111111111, 
10'b0000000001, 
10'b1111111110, 
10'b1111111110, 
10'b0000000001, 
10'b0000000110, 
10'b0000000011, 
10'b0000000101, 
10'b0000000001, 
10'b1111111011, 
10'b0000000001, 
10'b1111111011, 
10'b1111111101, 
10'b1111111100, 
10'b0000000000, 
10'b0000000000, 
10'b0000000010, 
10'b0000000001, 
10'b0000000010, 
10'b1111110110, 
10'b1111111011, 
10'b1111111111, 
10'b0000000000, 
10'b0000000111, 
10'b0000000111, 
10'b1111110111, 
10'b1111111110, 
10'b0000000100, 
10'b0000000110, 
10'b1111110111, 
10'b1111111011, 
10'b0000000000, 
10'b0000000100, 
10'b1111111101, 
10'b1111111101, 
10'b1111111110, 
10'b1111111111, 
10'b0000000110, 
10'b0000000101, 
10'b1111111111, 
10'b1111111101, 
10'b0000000100, 
10'b0000000010, 
10'b0000000100, 
10'b1111111111, 
10'b1111111100, 
10'b1111111110, 
10'b1111111111, 
10'b1111111001, 
10'b0000000001, 
10'b1111111001, 
10'b0000000011, 
10'b1111111111, 
10'b1111111111, 
10'b0000000100, 
10'b0000000000, 
10'b1111111111, 
10'b0000000010, 
10'b0000000010, 
10'b0000000001, 
10'b0000000000, 
10'b0000000011, 
10'b1111111011, 
10'b0000001000, 
10'b0000000011, 
10'b1111110111, 
10'b0000000000, 
10'b1111111001, 
10'b1111111000, 
10'b1111110110, 
10'b1111111110, 
10'b1111111101, 
10'b1111111100, 
10'b0000000010, 
10'b0000000000, 
10'b1111111001, 
10'b0000000001, 
10'b1111111100, 
10'b1111111100, 
10'b1111111101, 
10'b1111111101, 
10'b1111111100, 
10'b0000000000, 
10'b1111111110, 
10'b0000000100, 
10'b1111111100, 
10'b0000000001, 
10'b0000000000, 
10'b0000000010, 
10'b0000000110, 
10'b0000000000, 
10'b1111111011, 
10'b1111111101, 
10'b0000000011, 
10'b0000000100, 
10'b1111110101, 
10'b0000000010, 
10'b0000000000, 
10'b1111110111, 
10'b0000000101, 
10'b1111111101, 
10'b0000000000, 
10'b1111111011, 
10'b0000000101, 
10'b0000000011, 
10'b1111110100, 
10'b0000000100, 
10'b0000000010, 
10'b0000000010, 
10'b0000001001, 
10'b0000000010, 
10'b0000000101, 
10'b1111111011, 
10'b0000000001, 
10'b1111111110, 
10'b0000000010, 
10'b0000000111, 
10'b0000000011, 
10'b1111110101, 
10'b0000000101, 
10'b1111111101, 
10'b0000000001, 
10'b1111111011, 
10'b1111111010, 
10'b0000000001, 
10'b0000000011, 
10'b0000000001, 
10'b1111111110, 
10'b1111110110, 
10'b0000000010, 
10'b0000000000, 
10'b0000000100, 
10'b0000000000, 
10'b0000000001, 
10'b0000000100, 
10'b0000000100, 
10'b1111111101, 
10'b0000000011, 
10'b1111111011, 
10'b1111111011, 
10'b1111111101, 
10'b0000000101, 
10'b1111111100, 
10'b1111111010, 
10'b0000000000, 
10'b0000000011, 
10'b0000000100, 
10'b1111111100, 
10'b1111110111, 
10'b1111110111, 
10'b0000000011, 
10'b0000000000, 
10'b0000000101, 
10'b0000000100, 
10'b0000000011, 
10'b0000000101, 
10'b1111111101, 
10'b1111111111, 
10'b0000000001, 
10'b0000000010, 
10'b0000000100, 
10'b0000000101, 
10'b0000000110, 
10'b1111111011, 
10'b0000000000, 
10'b0000000110, 
10'b0000000100, 
10'b0000000100, 
10'b1111111111, 
10'b1111111010, 
10'b1111111110, 
10'b1111111110, 
10'b1111111011, 
10'b1111111000, 
10'b0000000100, 
10'b0000000011, 
10'b0000000101, 
10'b0000000000, 
10'b1111111100, 
10'b1111111110, 
10'b1111111100, 
10'b0000000000, 
10'b0000000000, 
10'b0000000101, 
10'b0000000010, 
10'b1111110111, 
10'b1111111011, 
10'b1111111010, 
10'b1111111111, 
10'b1111111000, 
10'b1111111110, 
10'b1111111101, 
10'b0000000001, 
10'b0000000000, 
10'b0000000001, 
10'b1111110110, 
10'b1111111111, 
10'b0000000100, 
10'b0000000110, 
10'b1111111111, 
10'b1111111000, 
10'b0000000011, 
10'b1111111110, 
10'b0000000101, 
10'b1111111111, 
10'b1111110110, 
10'b1111111101, 
10'b0000000000, 
10'b1111111000, 
10'b1111111111, 
10'b0000000101, 
10'b1111111101, 
10'b1111111111, 
10'b0000000101, 
10'b0000000001, 
10'b1111111101, 
10'b0000000101, 
10'b1111111101, 
10'b0000000010, 
10'b0000000000, 
10'b1111111001, 
10'b0000000101, 
10'b1111111100, 
10'b0000000000, 
10'b0000000000, 
10'b1111111101, 
10'b1111111110, 
10'b0000000011, 
10'b0000000000, 
10'b0000000001, 
10'b0000000010, 
10'b1111111100, 
10'b0000000001, 
10'b1111111010, 
10'b1111111111, 
10'b1111111100, 
10'b1111111100, 
10'b1111111011, 
10'b0000000000, 
10'b0000000010, 
10'b0000000001, 
10'b1111111101, 
10'b1111111011, 
10'b0000000101, 
10'b1111111100, 
10'b0000000000, 
10'b0000000110, 
10'b0000000000, 
10'b1111111001, 
10'b0000000100, 
10'b1111111011, 
10'b0000000010, 
10'b0000000001, 
10'b0000000010, 
10'b0000000100, 
10'b1111111011, 
10'b0000000001, 
10'b1111111100, 
10'b1111111010, 
10'b0000000011, 
10'b1111111001, 
10'b0000000101, 
10'b0000000001, 
10'b1111111101, 
10'b1111111001, 
10'b1111111101, 
10'b0000000101, 
10'b1111111100, 
10'b0000000000, 
10'b1111111101, 
10'b0000000110, 
10'b1111111110, 
10'b0000000000, 
10'b0000000011, 
10'b1111111100, 
10'b1111111100, 
10'b0000000001, 
10'b0000000000, 
10'b1111111000, 
10'b0000000110, 
10'b1111111110, 
10'b0000000110, 
10'b0000000011, 
10'b0000000011, 
10'b1111111011, 
10'b1111111110, 
10'b1111111110, 
10'b1111111101, 
10'b1111111111, 
10'b0000000011, 
10'b1111111100, 
10'b0000000011, 
10'b0000000000, 
10'b0000000001, 
10'b0000000011, 
10'b0000000101, 
10'b0000000010, 
10'b1111111100, 
10'b0000000001, 
10'b1111111000, 
10'b0000000010, 
10'b1111111101, 
10'b0000000011, 
10'b1111111101, 
10'b1111111100, 
10'b0000000010, 
10'b1111111011, 
10'b1111111100, 
10'b1111111010, 
10'b0000000000, 
10'b1111111100, 
10'b0000000111, 
10'b1111111111, 
10'b1111111100, 
10'b1111111111, 
10'b0000000010, 
10'b0000000010, 
10'b0000000101, 
10'b1111111101, 
10'b1111111010, 
10'b0000000000, 
10'b1111111011, 
10'b1111111101, 
10'b1111111001, 
10'b0000000011, 
10'b0000001000, 
10'b0000000011, 
10'b0000000101, 
10'b1111111111, 
10'b1111111100, 
10'b0000000100, 
10'b1111111110, 
10'b0000000101, 
10'b1111111101, 
10'b0000000001, 
10'b1111111010, 
10'b0000001000, 
10'b0000000111, 
10'b1111111100, 
10'b1111110101, 
10'b0000000000, 
10'b1111111011, 
10'b0000001000, 
10'b1111111111, 
10'b1111111100, 
10'b0000000000, 
10'b1111111100, 
10'b1111111100, 
10'b1111111101, 
10'b1111110110, 
10'b0000000000, 
10'b1111110110, 
10'b1111111101, 
10'b0000000000, 
10'b0000000010, 
10'b1111111100, 
10'b1111111111, 
10'b0000000001, 
10'b1111111101, 
10'b1111110101, 
10'b1111111101, 
10'b0000000001, 
10'b0000000001, 
10'b0000000010, 
10'b0000000010, 
10'b1111110111, 
10'b1111111101, 
10'b0000000101, 
10'b1111111001, 
10'b1111111101, 
10'b0000000111, 
10'b1111111100, 
10'b0000000000, 
10'b1111111100, 
10'b0000000001, 
10'b1111111110, 
10'b1111111101, 
10'b0000000101, 
10'b1111111001, 
10'b1111111101, 
10'b0000000100, 
10'b0000000101, 
10'b1111111110, 
10'b0000000010, 
10'b1111111110, 
10'b1111110111, 
10'b1111111101, 
10'b0000000001, 
10'b1111111100, 
10'b1111111111, 
10'b1111111110, 
10'b1111111100, 
10'b0000000100, 
10'b1111111100, 
10'b1111111100, 
10'b0000000000, 
10'b1111111110, 
10'b0000000010, 
10'b1111111010, 
10'b0000000101, 
10'b0000000011, 
10'b0000000000, 
10'b1111111111, 
10'b1111111011, 
10'b1111111010, 
10'b1111111100, 
10'b1111111101, 
10'b1111111110, 
10'b0000000001, 
10'b0000000111, 
10'b1111111101, 
10'b1111111000, 
10'b0000000111, 
10'b1111111100, 
10'b1111111111, 
10'b0000000001, 
10'b0000000011, 
10'b1111111011, 
10'b1111111100, 
10'b1111111110, 
10'b0000000011, 
10'b1111111100, 
10'b0000000011, 
10'b0000000011, 
10'b1111111010, 
10'b0000000000, 
10'b0000000000, 
10'b1111111110, 
10'b1111111101, 
10'b0000000000, 
10'b1111111110, 
10'b0000000001, 
10'b0000000001, 
10'b1111111010, 
10'b1111111100, 
10'b0000000000, 
10'b0000000011, 
10'b1111111001, 
10'b1111110111, 
10'b1111111100, 
10'b1111111110, 
10'b1111111110, 
10'b1111111111, 
10'b1111111011, 
10'b0000000010, 
10'b0000000010, 
10'b1111111100, 
10'b0000000011, 
10'b1111111111, 
10'b1111111101, 
10'b0000000101, 
10'b1111111100, 
10'b1111111110, 
10'b1111111100, 
10'b0000000001, 
10'b0000000100, 
10'b1111111111, 
10'b0000000010, 
10'b1111110110, 
10'b0000000000, 
10'b1111111100, 
10'b1111111101, 
10'b0000000100, 
10'b1111111010, 
10'b0000000010, 
10'b1111111101, 
10'b0000000000, 
10'b0000000000, 
10'b1111111001, 
10'b1111111111, 
10'b0000000000, 
10'b1111111011, 
10'b0000000001, 
10'b0000000101, 
10'b1111111100, 
10'b0000000011, 
10'b1111111110, 
10'b0000000110, 
10'b1111110101, 
10'b1111110101, 
10'b0000000011, 
10'b1111111101, 
10'b0000000001, 
10'b1111111011, 
10'b1111111110, 
10'b0000000011, 
10'b0000000001, 
10'b1111111111, 
10'b0000000001, 
10'b1111111100, 
10'b0000000100, 
10'b1111111111, 
10'b1111111100, 
10'b0000000010, 
10'b1111111111, 
10'b0000000000, 
10'b0000000011, 
10'b1111111001, 
10'b1111111100, 
10'b1111110101, 
10'b0000000010, 
10'b1111111001, 
10'b0000000011, 
10'b0000000010, 
10'b1111111111, 
10'b1111111011, 
10'b1111111100, 
10'b0000000011, 
10'b1111111111, 
10'b1111110111, 
10'b0000000110, 
10'b1111110111, 
10'b1111111011, 
10'b1111111111, 
10'b0000000000, 
10'b1111111010, 
10'b1111111101, 
10'b1111111111, 
10'b1111111111, 
10'b1111111110, 
10'b1111111111, 
10'b1111111100, 
10'b0000000111, 
10'b1111111110, 
10'b0000000000, 
10'b0000000000, 
10'b1111111110, 
10'b0000000001, 
10'b0000000000, 
10'b1111111110, 
10'b1111111110, 
10'b0000000001, 
10'b0000000000, 
10'b0000000001, 
10'b0000000010, 
10'b1111111011, 
10'b0000000111, 
10'b1111111101, 
10'b0000000001, 
10'b1111111101, 
10'b0000000010, 
10'b1111111010, 
10'b1111111011, 
10'b1111111000, 
10'b1111111110, 
10'b1111110101, 
10'b1111111111, 
10'b1111111100, 
10'b1111111010, 
10'b1111111011, 
10'b1111111101, 
10'b1111111100, 
10'b0000000101, 
10'b1111110101, 
10'b0000001000, 
10'b1111111110, 
10'b1111111011, 
10'b1111111110, 
10'b1111111001, 
10'b0000000001, 
10'b0000000010, 
10'b1111111010, 
10'b0000000001, 
10'b1111111000, 
10'b0000000100, 
10'b1111111001, 
10'b0000000001, 
10'b1111111101, 
10'b1111111110, 
10'b0000000101, 
10'b0000000100, 
10'b1111111100, 
10'b0000000100, 
10'b0000000001, 
10'b0000000001, 
10'b0000000110, 
10'b0000000011, 
10'b1111111100, 
10'b1111111100, 
10'b0000000101, 
10'b0000000101, 
10'b0000000000, 
10'b0000000011, 
10'b0000000001, 
10'b0000000001, 
10'b1111111110, 
10'b0000000100, 
10'b1111111111, 
10'b0000000000, 
10'b0000000001, 
10'b0000001001, 
10'b1111111010, 
10'b1111111101, 
10'b0000000000, 
10'b0000000100, 
10'b0000000100, 
10'b1111111011, 
10'b1111111010, 
10'b0000000000, 
10'b0000000001, 
10'b0000000000, 
10'b0000000001, 
10'b0000000010, 
10'b0000000001, 
10'b0000000100, 
10'b1111111111, 
10'b0000000000, 
10'b0000000100, 
10'b1111111111, 
10'b1111111110, 
10'b0000000001, 
10'b1111111001, 
10'b0000000000, 
10'b0000000010, 
10'b1111111010, 
10'b0000000111, 
10'b1111111111, 
10'b0000000001, 
10'b1111111111, 
10'b1111111110, 
10'b1111111110, 
10'b0000000011, 
10'b0000000111, 
10'b0000000000, 
10'b0000000011, 
10'b0000001000, 
10'b1111111001, 
10'b0000000011, 
10'b0000000100, 
10'b1111111011, 
10'b0000000000, 
10'b0000000100, 
10'b0000000000, 
10'b0000000011, 
10'b1111111111, 
10'b0000000110, 
10'b0000000010, 
10'b1111111101, 
10'b1111111000, 
10'b1111111011, 
10'b0000000001, 
10'b0000000000, 
10'b1111111111, 
10'b0000000010, 
10'b0000000010, 
10'b0000000010, 
10'b1111111000, 
10'b0000000001, 
10'b0000000011, 
10'b1111111001, 
10'b1111111100, 
10'b1111111110, 
10'b0000000110, 
10'b0000000110, 
10'b1111111111, 
10'b0000000011, 
10'b1111111001, 
10'b1111111101, 
10'b1111111101, 
10'b1111111111, 
10'b0000000000, 
10'b1111110111, 
10'b0000000011, 
10'b1111111110, 
10'b1111111110, 
10'b1111111010, 
10'b0000000000, 
10'b1111111111, 
10'b0000001001, 
10'b1111111000, 
10'b0000000010, 
10'b0000000000, 
10'b1111111100, 
10'b1111111101, 
10'b0000000001, 
10'b1111111010, 
10'b1111111100, 
10'b1111111000, 
10'b1111111110, 
10'b0000000011, 
10'b0000000110, 
10'b1111111011, 
10'b1111111110, 
10'b0000000001, 
10'b0000000101, 
10'b1111111101, 
10'b1111111111, 
10'b1111111111, 
10'b0000000101, 
10'b1111110111, 
10'b0000000101, 
10'b1111111100, 
10'b1111110111, 
10'b1111111011, 
10'b0000001000, 
10'b1111111001, 
10'b1111111110, 
10'b1111111000, 
10'b0000000011, 
10'b0000000111, 
10'b0000000111, 
10'b1111111011, 
10'b0000000000, 
10'b1111110111, 
10'b0000000011, 
10'b1111111100, 
10'b0000000100, 
10'b0000000000, 
10'b0000000010, 
10'b1111111100, 
10'b1111111100, 
10'b1111111011, 
10'b0000000001, 
10'b0000000010, 
10'b0000000110, 
10'b0000000001, 
10'b1111111100, 
10'b1111111110, 
10'b1111111001, 
10'b0000000101, 
10'b0000000011, 
10'b1111111010, 
10'b1111111110, 
10'b1111110111, 
10'b0000000101, 
10'b1111111001, 
10'b0000000110, 
10'b1111111011, 
10'b0000000001, 
10'b0000000000, 
10'b0000000101, 
10'b1111111011, 
10'b1111111010, 
10'b0000000101, 
10'b1111111100, 
10'b0000000000, 
10'b1111111010, 
10'b0000000000, 
10'b1111111101, 
10'b0000000011, 
10'b1111111101, 
10'b1111111100, 
10'b1111111101, 
10'b0000000011, 
10'b1111111101, 
10'b1111111110, 
10'b0000000010, 
10'b0000000100, 
10'b1111111000, 
10'b0000000000, 
10'b0000000000, 
10'b1111110111, 
10'b1111111110, 
10'b0000000110, 
10'b0000000011, 
10'b1111111000, 
10'b0000000011, 
10'b1111110010, 
10'b1111111001, 
10'b1111111010, 
10'b0000000000, 
10'b1111110111, 
10'b1111111101, 
10'b0000000000, 
10'b1111111101, 
10'b0000000111, 
10'b0000000001, 
10'b0000000000, 
10'b0000000000, 
10'b0000001001, 
10'b1111111010, 
10'b1111111010, 
10'b0000000001, 
10'b0000000101, 
10'b0000000100, 
10'b0000000100, 
10'b1111111100, 
10'b1111111010, 
10'b0000000000, 
10'b1111111011, 
10'b0000000001, 
10'b0000000001, 
10'b0000000000, 
10'b1111111000, 
10'b1111111000, 
10'b1111111111, 
10'b1111111110, 
10'b1111111110, 
10'b1111111000, 
10'b0000000001, 
10'b1111111101, 
10'b1111110110, 
10'b1111111011, 
10'b0000000101, 
10'b1111111001, 
10'b0000000100, 
10'b0000001000, 
10'b0000000111, 
10'b1111111111, 
10'b1111111010, 
10'b0000000011, 
10'b1111111010, 
10'b1111111101, 
10'b0000000011, 
10'b1111111111, 
10'b1111111110, 
10'b1111111110, 
10'b0000000100

};
localparam logic signed [9:0] dlBiases [9:0] = {
10'b0000000101, 
10'b1111111111, 
10'b1111111111, 
10'b1111111110, 
10'b1111111110, 
10'b1111111111, 
10'b1111111111, 
10'b0000000010, 
10'b1111111010, 
10'b1111111111 

};
localparam logic signed [9:0] convWeights [0:17] = {
10'b0000000011, 
10'b0000001111, 
10'b1111111000, 
10'b0000000010, 
10'b0000000000, 
10'b0000010000, 
10'b0000001100, 
10'b0000000110, 
10'b1111111000, 
10'b0000001011, 
10'b1111111101, 
10'b0000000110, 
10'b0000001111, 
10'b0000000101, 
10'b0000001100, 
10'b1111111111, 
10'b0000000101, 
10'b0000000011

};
localparam logic signed [9:0] convBiases [1:0] = {
10'b0000000000, 
10'b0000000000

};
endpackage