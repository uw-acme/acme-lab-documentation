package data22_11;
localparam logic signed [21:0] dlWeights [0:1279] = {
22'b0000000000001000001110, 
22'b0000000000000000010100, 
22'b1111111111111001110000, 
22'b0000000000000000001101, 
22'b1111111111111101111010, 
22'b0000000000000100010010, 
22'b0000000000000010000001, 
22'b1111111111111001101000, 
22'b0000000000000001011101, 
22'b0000000000000101010111, 
22'b0000000000000101011000, 
22'b1111111111110111101111, 
22'b1111111111110011110111, 
22'b1111111111111010100110, 
22'b0000000000000011000100, 
22'b1111111111111100001001, 
22'b1111111111111101100110, 
22'b1111111111111111000010, 
22'b1111111111111110011000, 
22'b1111111111111111111001, 
22'b0000000000000011110110, 
22'b1111111111111000010110, 
22'b0000000000000001101110, 
22'b0000000000000010100100, 
22'b1111111111111110111101, 
22'b0000000000000000001010, 
22'b1111111111111101111001, 
22'b0000000000000001000111, 
22'b0000000000000010000101, 
22'b0000000000001000000110, 
22'b0000000000010010010110, 
22'b1111111111110010010101, 
22'b1111111111111000001100, 
22'b1111111111110110101000, 
22'b1111111111111000100011, 
22'b0000000000000011111001, 
22'b1111111111111111001010, 
22'b0000000000000101001101, 
22'b1111111111111101101111, 
22'b0000000000000110100100, 
22'b0000000000000100111111, 
22'b1111111111111011101011, 
22'b1111111111111111011101, 
22'b1111111111111010100101, 
22'b0000000000000000001011, 
22'b1111111111111100111101, 
22'b0000000000000101100101, 
22'b1111111111111011001101, 
22'b1111111111111100011011, 
22'b0000000000000000010100, 
22'b0000000000001011101011, 
22'b1111111111111011011010, 
22'b1111111111110111110001, 
22'b1111111111110101010011, 
22'b1111111111111010110100, 
22'b0000000000000011000110, 
22'b1111111111111111010010, 
22'b0000000000000100000100, 
22'b0000000000000010000011, 
22'b0000000000000011010010, 
22'b0000000000000111110001, 
22'b1111111111111001101010, 
22'b0000000000000010000110, 
22'b0000000000000010001001, 
22'b1111111111111010100101, 
22'b0000000000000111010010, 
22'b0000000000000110110100, 
22'b0000000000000000000101, 
22'b0000000000000101100110, 
22'b1111111111111101011100, 
22'b0000000000000000000111, 
22'b0000000000000110101101, 
22'b1111111111111000111111, 
22'b1111111111111011000111, 
22'b1111111111111010111010, 
22'b0000000000000011001011, 
22'b1111111111111110101110, 
22'b0000000000000101101000, 
22'b1111111111111000100010, 
22'b1111111111111010001111, 
22'b1111111111111101100101, 
22'b1111111111111100101001, 
22'b1111111111111000110001, 
22'b0000000000000011010111, 
22'b1111111111111011101100, 
22'b0000000000000100010001, 
22'b0000000000000000000000, 
22'b1111111111111010100111, 
22'b1111111111111110001111, 
22'b1111111111111100011101, 
22'b0000000000000001001000, 
22'b0000000000000000100010, 
22'b1111111111111100100110, 
22'b0000000000000000111000, 
22'b1111111111110111000001, 
22'b1111111111111110010110, 
22'b1111111111111000010110, 
22'b0000000000001010000010, 
22'b1111111111110111101101, 
22'b1111111111110110010100, 
22'b0000000000000000101010, 
22'b0000000000001001100001, 
22'b0000000000000000001010, 
22'b0000000000000001000110, 
22'b1111111111111011001101, 
22'b1111111111111111001110, 
22'b1111111111111010010011, 
22'b1111111111111010101001, 
22'b0000000000000011011110, 
22'b1111111111111001110000, 
22'b0000000000000000111001, 
22'b0000000000000101010100, 
22'b0000000000000001000111, 
22'b0000000000000100000101, 
22'b1111111111111000000100, 
22'b1111111111111100110011, 
22'b1111111111110111100100, 
22'b0000000000000011100011, 
22'b1111111111111010101111, 
22'b0000000000000010000011, 
22'b1111111111111010000011, 
22'b1111111111111110001110, 
22'b0000000000000000100011, 
22'b0000000000000010011010, 
22'b1111111111111000011101, 
22'b1111111111111101111010, 
22'b1111111111111000100100, 
22'b1111111111111100110001, 
22'b0000000000000000000100, 
22'b0000000000000010101001, 
22'b1111111111111010110101, 
22'b1111111111111101111101, 
22'b1111111111111100101010, 
22'b0000000000001000111101, 
22'b1111111111111010011010, 
22'b1111111111110101110001, 
22'b1111111111111011010010, 
22'b0000000000001010001001, 
22'b1111111111111110010011, 
22'b0000000000000001100000, 
22'b1111111111111111100110, 
22'b1111111111111101011110, 
22'b0000000000000000011111, 
22'b0000000000000001100000, 
22'b0000000000000110011111, 
22'b1111111111111110101100, 
22'b1111111111110111100100, 
22'b0000000000000110100111, 
22'b1111111111111110010000, 
22'b0000000000000010001100, 
22'b0000000000000000101001, 
22'b0000000000000010101011, 
22'b0000000000000100101010, 
22'b1111111111111111101011, 
22'b0000000000000010100111, 
22'b1111111111111011010101, 
22'b1111111111100111111110, 
22'b0000000000000110011001, 
22'b1111111111111110100100, 
22'b0000000000000011001100, 
22'b0000000000000101000110, 
22'b1111111111111110001000, 
22'b1111111111110111101111, 
22'b0000000000000101111011, 
22'b0000000000000110111001, 
22'b1111111111111100100110, 
22'b0000000000001000000101, 
22'b1111111111111110001011, 
22'b0000000000000001010111, 
22'b1111111111111111011001, 
22'b0000000000000100101110, 
22'b1111111111111111100000, 
22'b1111111111111110001001, 
22'b1111111111110101000101, 
22'b0000000000000000100110, 
22'b0000000000000001110011, 
22'b1111111111111101010111, 
22'b1111111111111111001000, 
22'b1111111111111100011010, 
22'b0000000000000100101100, 
22'b0000000000000111100001, 
22'b1111111111111000100001, 
22'b1111111111111111011100, 
22'b1111111111111101000101, 
22'b0000000000000111100101, 
22'b1111111111111111101101, 
22'b0000000000000100011100, 
22'b1111111111111100011111, 
22'b0000000000000110010111, 
22'b0000000000000000001111, 
22'b0000000000000111100001, 
22'b1111111111110100111000, 
22'b1111111111111011010110, 
22'b1111111111110111100011, 
22'b1111111111111111110010, 
22'b0000000000000010111011, 
22'b0000000000000001010110, 
22'b0000000000000011010100, 
22'b0000000000000100111111, 
22'b1111111111111110100100, 
22'b0000000000000110100011, 
22'b1111111111110111101000, 
22'b1111111111111100100100, 
22'b1111111111111011101001, 
22'b1111111111111111111100, 
22'b0000000000000000010110, 
22'b0000000000000000000111, 
22'b1111111111111110111110, 
22'b0000000000000000101011, 
22'b1111111111111100110000, 
22'b1111111111111110001011, 
22'b1111111111111110101010, 
22'b1111111111111110100101, 
22'b1111111111111001011001, 
22'b1111111111111111100001, 
22'b0000000000000000110101, 
22'b0000000000000110101000, 
22'b1111111111111101000100, 
22'b0000000000000000011111, 
22'b0000000000000001011011, 
22'b1111111111111011101111, 
22'b1111111111111110011001, 
22'b1111111111111001110110, 
22'b0000000000000101111100, 
22'b1111111111111001101110, 
22'b0000000000000111101011, 
22'b1111111111111010010011, 
22'b0000000000000000100111, 
22'b1111111111111101010110, 
22'b1111111111110111011110, 
22'b0000000000000101000100, 
22'b0000000000000111010110, 
22'b1111111111111001111111, 
22'b0000000000000010001111, 
22'b1111111111111111010000, 
22'b0000000000000000011101, 
22'b1111111111111100101001, 
22'b0000000000000101000100, 
22'b0000000000000001111110, 
22'b0000000000000001100111, 
22'b0000000000000000000110, 
22'b1111111111111100101001, 
22'b0000000000000010101001, 
22'b0000000000000011110111, 
22'b0000000000000010100001, 
22'b1111111111111101011001, 
22'b1111111111111010101100, 
22'b1111111111111101111101, 
22'b0000000000000011110010, 
22'b1111111111111011010010, 
22'b0000000000000010011001, 
22'b0000000000000010001101, 
22'b1111111111111101100111, 
22'b1111111111111011111111, 
22'b1111111111110111101000, 
22'b1111111111111100101100, 
22'b0000000000000000010101, 
22'b0000000000000000000010, 
22'b1111111111110110010101, 
22'b1111111111111001011110, 
22'b1111111111111000000000, 
22'b0000000000000001011000, 
22'b0000000000000000111111, 
22'b0000000000000010110101, 
22'b1111111111110101010110, 
22'b0000000000000000101110, 
22'b0000000000000011100011, 
22'b1111111111111001011100, 
22'b0000000000000000010011, 
22'b1111111111111111001110, 
22'b0000000000000000111100, 
22'b0000000000000101111000, 
22'b0000000000000001101000, 
22'b0000000000000000111011, 
22'b1111111111111110111000, 
22'b1111111111111001100010, 
22'b1111111111111000111000, 
22'b0000000000001000011110, 
22'b1111111111110111001011, 
22'b0000000000000000101010, 
22'b1111111111111111101000, 
22'b0000000000000000010000, 
22'b0000000000000010110101, 
22'b1111111111111110010100, 
22'b0000000000000001000110, 
22'b1111111111111100100001, 
22'b0000000000000011010000, 
22'b1111111111111111111101, 
22'b0000000000000100100011, 
22'b0000000000000010111011, 
22'b1111111111111100100010, 
22'b0000000000000011101101, 
22'b0000000000000011101110, 
22'b0000000000000000001011, 
22'b0000000000000010110100, 
22'b1111111111111100111101, 
22'b1111111111110110010000, 
22'b1111111111111111011011, 
22'b1111111111111010100010, 
22'b1111111111111101110101, 
22'b0000000000000001001101, 
22'b0000000000000110011001, 
22'b0000000000000001100001, 
22'b0000000000000010111100, 
22'b1111111111111101110000, 
22'b0000000000000001010000, 
22'b0000000000000010101011, 
22'b1111111111111101111000, 
22'b0000000000000011001100, 
22'b0000000000000110011100, 
22'b0000000000000011111111, 
22'b0000000000000010011000, 
22'b1111111111111110110011, 
22'b0000000000000001100000, 
22'b0000000000000100101110, 
22'b0000000000000010101001, 
22'b1111111111111000011010, 
22'b0000000000000000100101, 
22'b1111111111111110101000, 
22'b1111111111111111110110, 
22'b0000000000000100001011, 
22'b1111111111110111011011, 
22'b1111111111111011100110, 
22'b0000000000000011011000, 
22'b0000000000000110111000, 
22'b0000000000000000100110, 
22'b0000000000000110111111, 
22'b1111111111110111110010, 
22'b0000000000000000010000, 
22'b0000000000000011110101, 
22'b0000000000001000111011, 
22'b1111111111110111100010, 
22'b1111111111111101010000, 
22'b1111111111110101110110, 
22'b1111111111111110000001, 
22'b0000000000000011001111, 
22'b1111111111111011111110, 
22'b0000000000000001011000, 
22'b1111111111111101001110, 
22'b1111111111111011010000, 
22'b0000000000000011110001, 
22'b1111111111111101010000, 
22'b1111111111111110011100, 
22'b1111111111111010000010, 
22'b0000000000000001001111, 
22'b1111111111111101110010, 
22'b0000000000000001111010, 
22'b1111111111111100101100, 
22'b0000000000000101000110, 
22'b1111111111111011100111, 
22'b0000000000000101000111, 
22'b1111111111111101101010, 
22'b1111111111110100110101, 
22'b0000000000000001100110, 
22'b0000000000000100110101, 
22'b0000000000000000010110, 
22'b0000000000000000110110, 
22'b0000000000000001000010, 
22'b0000000000000101001010, 
22'b1111111111111100111000, 
22'b0000000000000001011111, 
22'b1111111111111000001111, 
22'b0000000000000100000010, 
22'b0000000000000100100010, 
22'b0000000000000000100111, 
22'b1111111111111101111000, 
22'b0000000000000010100111, 
22'b1111111111111110000101, 
22'b0000000000000010001010, 
22'b0000000000000001000111, 
22'b0000000000000000000010, 
22'b0000000000000000110000, 
22'b1111111111111011001110, 
22'b0000000000000001100000, 
22'b1111111111111110100111, 
22'b0000000000000001001111, 
22'b0000000000000110101001, 
22'b0000000000000100010110, 
22'b1111111111111111010010, 
22'b1111111111111001101010, 
22'b0000000000000011100100, 
22'b1111111111111000101010, 
22'b1111111111111101111111, 
22'b1111111111111100111101, 
22'b1111111111111111110111, 
22'b0000000000000101011110, 
22'b1111111111111110010110, 
22'b0000000000000000000101, 
22'b0000000000000111110000, 
22'b1111111111111110100010, 
22'b1111111111111110100010, 
22'b1111111111111101111001, 
22'b1111111111111111011000, 
22'b0000000000000100001001, 
22'b1111111111111010010000, 
22'b1111111111111101001111, 
22'b1111111111111101010101, 
22'b1111111111111001110101, 
22'b1111111111111011110001, 
22'b1111111111110111101001, 
22'b1111111111111100101101, 
22'b1111111111111100111001, 
22'b1111111111110111111110, 
22'b0000000000000110001100, 
22'b1111111111111001111111, 
22'b0000000000000010001100, 
22'b1111111111111010101111, 
22'b1111111111111010110010, 
22'b0000000000000011110111, 
22'b0000000000000000000111, 
22'b1111111111111010010100, 
22'b0000000000000001011101, 
22'b1111111111111001011100, 
22'b0000000000000101001001, 
22'b0000000000000010010001, 
22'b1111111111111101101000, 
22'b1111111111111011110111, 
22'b1111111111111100000110, 
22'b0000000000000011001110, 
22'b1111111111111010000000, 
22'b0000000000000000010101, 
22'b0000000000000101001001, 
22'b0000000000000010110000, 
22'b0000000000000011011010, 
22'b1111111111111010011001, 
22'b0000000000000110011110, 
22'b0000000000000100111011, 
22'b0000000000000000110010, 
22'b0000000000000111010000, 
22'b0000000000000000111010, 
22'b1111111111110111001111, 
22'b0000000000000110110000, 
22'b0000000000000010100111, 
22'b0000000000000101100110, 
22'b1111111111111000111000, 
22'b1111111111111110100111, 
22'b0000000000000001110011, 
22'b1111111111111010011101, 
22'b1111111111111011001001, 
22'b1111111111111011011100, 
22'b1111111111111100101110, 
22'b0000000000000111010100, 
22'b0000000000000000011011, 
22'b0000000000000011010001, 
22'b0000000000000000011001, 
22'b0000000000000110000101, 
22'b0000000000000101110001, 
22'b1111111111111000011111, 
22'b1111111111111010110000, 
22'b0000000000000100011010, 
22'b1111111111111011110111, 
22'b1111111111111110110000, 
22'b1111111111111110110001, 
22'b0000000000000100000111, 
22'b0000000000000001100011, 
22'b1111111111111111101110, 
22'b1111111111111010101011, 
22'b0000000000000100111101, 
22'b1111111111111110010101, 
22'b0000000000000101011100, 
22'b0000000000000001111010, 
22'b0000000000000010101010, 
22'b1111111111111101111100, 
22'b0000000000000000100011, 
22'b0000000000000101011100, 
22'b1111111111111110111011, 
22'b1111111111111111101000, 
22'b1111111111111111010001, 
22'b1111111111111011001111, 
22'b0000000000001000000010, 
22'b0000000000000001001101, 
22'b1111111111111100001011, 
22'b1111111111111111010101, 
22'b0000000000000001110001, 
22'b1111111111111110100111, 
22'b1111111111111110100010, 
22'b0000000000000001001000, 
22'b0000000000000110010110, 
22'b0000000000000011100011, 
22'b0000000000000101101100, 
22'b0000000000000001111110, 
22'b1111111111111011010000, 
22'b0000000000000001010000, 
22'b1111111111111011010001, 
22'b1111111111111101010100, 
22'b1111111111111100001001, 
22'b0000000000000000000010, 
22'b0000000000000000101100, 
22'b0000000000000010101110, 
22'b0000000000000001100111, 
22'b0000000000000010000010, 
22'b1111111111110110011100, 
22'b1111111111111011000000, 
22'b1111111111111111000011, 
22'b0000000000000000111000, 
22'b0000000000000111101101, 
22'b0000000000000111100011, 
22'b1111111111110111100110, 
22'b1111111111111110111111, 
22'b0000000000000100001001, 
22'b0000000000000110101100, 
22'b1111111111110111100110, 
22'b1111111111111011010010, 
22'b0000000000000000111000, 
22'b0000000000000100101101, 
22'b1111111111111101000110, 
22'b1111111111111101110110, 
22'b1111111111111110010011, 
22'b1111111111111111101011, 
22'b0000000000000110101101, 
22'b0000000000000101010011, 
22'b1111111111111111011011, 
22'b1111111111111101101100, 
22'b0000000000000100101100, 
22'b0000000000000010010001, 
22'b0000000000000100010101, 
22'b1111111111111111001111, 
22'b1111111111111100001111, 
22'b1111111111111110001100, 
22'b1111111111111111001000, 
22'b1111111111111001010000, 
22'b0000000000000001011011, 
22'b1111111111111001100001, 
22'b0000000000000011001111, 
22'b1111111111111111000011, 
22'b1111111111111111001010, 
22'b0000000000000100000110, 
22'b0000000000000000100111, 
22'b1111111111111111010110, 
22'b0000000000000010101101, 
22'b0000000000000010000110, 
22'b0000000000000001101111, 
22'b0000000000000000110111, 
22'b0000000000000011000000, 
22'b1111111111111011111010, 
22'b0000000000001000000101, 
22'b0000000000000011111101, 
22'b1111111111110111010011, 
22'b0000000000000000100101, 
22'b1111111111111001000011, 
22'b1111111111111000110000, 
22'b1111111111110110101111, 
22'b1111111111111110010100, 
22'b1111111111111101010110, 
22'b1111111111111100000111, 
22'b0000000000000010110110, 
22'b0000000000000000100000, 
22'b1111111111111001111101, 
22'b0000000000000001010010, 
22'b1111111111111100001101, 
22'b1111111111111100100001, 
22'b1111111111111101000000, 
22'b1111111111111101111011, 
22'b1111111111111100110001, 
22'b0000000000000000100010, 
22'b1111111111111110010011, 
22'b0000000000000100101100, 
22'b1111111111111100000010, 
22'b0000000000000001101100, 
22'b0000000000000000110011, 
22'b0000000000000010110010, 
22'b0000000000000110110011, 
22'b0000000000000000000011, 
22'b1111111111111011101010, 
22'b1111111111111101000001, 
22'b0000000000000011100101, 
22'b0000000000000100011101, 
22'b1111111111110101111010, 
22'b0000000000000010011011, 
22'b0000000000000000100111, 
22'b1111111111110111010100, 
22'b0000000000000101101011, 
22'b1111111111111101100010, 
22'b0000000000000000001001, 
22'b1111111111111011011100, 
22'b0000000000000101100001, 
22'b0000000000000011111001, 
22'b1111111111110100110101, 
22'b0000000000000100011100, 
22'b0000000000000010111111, 
22'b0000000000000010110010, 
22'b0000000000001001010011, 
22'b0000000000000010100111, 
22'b0000000000000101000101, 
22'b1111111111111011000110, 
22'b0000000000000001001001, 
22'b1111111111111110001001, 
22'b0000000000000010001001, 
22'b0000000000000111011000, 
22'b0000000000000011101101, 
22'b1111111111110101110100, 
22'b0000000000000101001101, 
22'b1111111111111101101100, 
22'b0000000000000001011011, 
22'b1111111111111011111010, 
22'b1111111111111010010010, 
22'b0000000000000001000110, 
22'b0000000000000011110001, 
22'b0000000000000001111011, 
22'b1111111111111110001100, 
22'b1111111111110110110001, 
22'b0000000000000010010100, 
22'b0000000000000000110111, 
22'b0000000000000100101000, 
22'b0000000000000000001100, 
22'b0000000000000001000101, 
22'b0000000000000100111010, 
22'b0000000000000100010001, 
22'b1111111111111101101101, 
22'b0000000000000011011100, 
22'b1111111111111011111011, 
22'b1111111111111011111101, 
22'b1111111111111101010001, 
22'b0000000000000101100100, 
22'b1111111111111100001110, 
22'b1111111111111010011111, 
22'b0000000000000000111011, 
22'b0000000000000011011110, 
22'b0000000000000100010010, 
22'b1111111111111100111010, 
22'b1111111111110111011100, 
22'b1111111111110111001110, 
22'b0000000000000011110100, 
22'b0000000000000000011111, 
22'b0000000000000101011100, 
22'b0000000000000100011011, 
22'b0000000000000011101110, 
22'b0000000000000101110000, 
22'b1111111111111101001110, 
22'b1111111111111111100000, 
22'b0000000000000001011011, 
22'b0000000000000010010101, 
22'b0000000000000100111001, 
22'b0000000000000101011100, 
22'b0000000000000110100001, 
22'b1111111111111011110011, 
22'b0000000000000000000010, 
22'b0000000000000110101001, 
22'b0000000000000100110111, 
22'b0000000000000100100010, 
22'b1111111111111111100111, 
22'b1111111111111010111111, 
22'b1111111111111110101000, 
22'b1111111111111110110100, 
22'b1111111111111011110001, 
22'b1111111111111000001000, 
22'b0000000000000100001111, 
22'b0000000000000011110000, 
22'b0000000000000101000011, 
22'b0000000000000000000100, 
22'b1111111111111100111101, 
22'b1111111111111110101110, 
22'b1111111111111100001101, 
22'b0000000000000000111101, 
22'b0000000000000000000101, 
22'b0000000000000101111010, 
22'b0000000000000010100110, 
22'b1111111111110111000101, 
22'b1111111111111011011100, 
22'b1111111111111010010110, 
22'b1111111111111111110010, 
22'b1111111111111000110000, 
22'b1111111111111110011110, 
22'b1111111111111101101000, 
22'b0000000000000001101111, 
22'b0000000000000000010011, 
22'b0000000000000001000111, 
22'b1111111111110110011011, 
22'b1111111111111111101000, 
22'b0000000000000100010100, 
22'b0000000000000110110001, 
22'b1111111111111111010101, 
22'b1111111111111000011111, 
22'b0000000000000011110011, 
22'b1111111111111110001100, 
22'b0000000000000101101010, 
22'b1111111111111111110100, 
22'b1111111111110110111111, 
22'b1111111111111101000011, 
22'b0000000000000000101100, 
22'b1111111111111000100111, 
22'b1111111111111111010101, 
22'b0000000000000101101001, 
22'b1111111111111101101000, 
22'b1111111111111111101011, 
22'b0000000000000101011111, 
22'b0000000000000001110110, 
22'b1111111111111101101110, 
22'b0000000000000101110001, 
22'b1111111111111101110001, 
22'b0000000000000010011001, 
22'b0000000000000000011011, 
22'b1111111111111001110100, 
22'b0000000000000101000010, 
22'b1111111111111100110110, 
22'b0000000000000000010011, 
22'b0000000000000000101001, 
22'b1111111111111101001111, 
22'b1111111111111110011001, 
22'b0000000000000011100010, 
22'b0000000000000000000100, 
22'b0000000000000001011010, 
22'b0000000000000010011010, 
22'b1111111111111100011101, 
22'b0000000000000001110101, 
22'b1111111111111010101101, 
22'b1111111111111111110111, 
22'b1111111111111100110110, 
22'b1111111111111100101000, 
22'b1111111111111011001001, 
22'b0000000000000000110000, 
22'b0000000000000010101000, 
22'b0000000000000001011110, 
22'b1111111111111101100001, 
22'b1111111111111011010100, 
22'b0000000000000101010011, 
22'b1111111111111100111110, 
22'b0000000000000000000010, 
22'b0000000000000110011110, 
22'b0000000000000000001000, 
22'b1111111111111001100101, 
22'b0000000000000100011010, 
22'b1111111111111011100110, 
22'b0000000000000010111011, 
22'b0000000000000001111110, 
22'b0000000000000010000010, 
22'b0000000000000100001110, 
22'b1111111111111011000011, 
22'b0000000000000001100101, 
22'b1111111111111100110001, 
22'b1111111111111010001011, 
22'b0000000000000011011100, 
22'b1111111111111001110101, 
22'b0000000000000101101011, 
22'b0000000000000001000101, 
22'b1111111111111101110000, 
22'b1111111111111001100100, 
22'b1111111111111101001111, 
22'b0000000000000101010011, 
22'b1111111111111100000110, 
22'b0000000000000000010100, 
22'b1111111111111101010010, 
22'b0000000000000110000001, 
22'b1111111111111110111100, 
22'b0000000000000000100110, 
22'b0000000000000011000010, 
22'b1111111111111100110101, 
22'b1111111111111100011000, 
22'b0000000000000001100000, 
22'b0000000000000000110011, 
22'b1111111111111000101000, 
22'b0000000000000110110100, 
22'b1111111111111110100101, 
22'b0000000000000110010100, 
22'b0000000000000011100010, 
22'b0000000000000011001001, 
22'b1111111111111011100001, 
22'b1111111111111110100001, 
22'b1111111111111110100000, 
22'b1111111111111101110000, 
22'b1111111111111111010110, 
22'b0000000000000011100010, 
22'b1111111111111100000111, 
22'b0000000000000011001100, 
22'b0000000000000000101110, 
22'b0000000000000001000101, 
22'b0000000000000011010011, 
22'b0000000000000101000010, 
22'b0000000000000010101010, 
22'b1111111111111100010000, 
22'b0000000000000001110101, 
22'b1111111111111000011111, 
22'b0000000000000010001001, 
22'b1111111111111101101000, 
22'b0000000000000011000101, 
22'b1111111111111101001001, 
22'b1111111111111100100111, 
22'b0000000000000010101010, 
22'b1111111111111011000110, 
22'b1111111111111100111111, 
22'b1111111111111010100110, 
22'b0000000000000000111011, 
22'b1111111111111100011010, 
22'b0000000000000111001101, 
22'b1111111111111111010011, 
22'b1111111111111100010001, 
22'b1111111111111111111000, 
22'b0000000000000010100100, 
22'b0000000000000010100001, 
22'b0000000000000101011111, 
22'b1111111111111101011111, 
22'b1111111111111010000000, 
22'b0000000000000000011010, 
22'b1111111111111011110110, 
22'b1111111111111101011100, 
22'b1111111111111001000000, 
22'b0000000000000011011000, 
22'b0000000000001000011010, 
22'b0000000000000011001110, 
22'b0000000000000101001110, 
22'b1111111111111111110010, 
22'b1111111111111100011001, 
22'b0000000000000100100000, 
22'b1111111111111110000111, 
22'b0000000000000101000110, 
22'b1111111111111101100110, 
22'b0000000000000001011101, 
22'b1111111111111010001100, 
22'b0000000000001000110001, 
22'b0000000000000111100100, 
22'b1111111111111100100111, 
22'b1111111111110101110011, 
22'b0000000000000000101110, 
22'b1111111111111011000110, 
22'b0000000000001000000111, 
22'b1111111111111111000001, 
22'b1111111111111100110110, 
22'b0000000000000000110101, 
22'b1111111111111100011000, 
22'b1111111111111100101011, 
22'b1111111111111101110110, 
22'b1111111111110110011111, 
22'b0000000000000000111100, 
22'b1111111111110110101001, 
22'b1111111111111101010101, 
22'b0000000000000000110110, 
22'b0000000000000010111010, 
22'b1111111111111100011110, 
22'b1111111111111111011100, 
22'b0000000000000001010000, 
22'b1111111111111101101101, 
22'b1111111111110101010001, 
22'b1111111111111101101011, 
22'b0000000000000001101010, 
22'b0000000000000001001011, 
22'b0000000000000010010101, 
22'b0000000000000010100010, 
22'b1111111111110111011100, 
22'b1111111111111101000001, 
22'b0000000000000101100011, 
22'b1111111111111001110011, 
22'b1111111111111101110001, 
22'b0000000000000111011101, 
22'b1111111111111100110001, 
22'b0000000000000000001101, 
22'b1111111111111100111001, 
22'b0000000000000001000010, 
22'b1111111111111110101111, 
22'b1111111111111101110011, 
22'b0000000000000101111100, 
22'b1111111111111001111110, 
22'b1111111111111101110011, 
22'b0000000000000100100101, 
22'b0000000000000101110100, 
22'b1111111111111110010101, 
22'b0000000000000010000101, 
22'b1111111111111110110000, 
22'b1111111111110111010001, 
22'b1111111111111101111000, 
22'b0000000000000001001001, 
22'b1111111111111100111000, 
22'b1111111111111111110000, 
22'b1111111111111110000000, 
22'b1111111111111100111001, 
22'b0000000000000100110101, 
22'b1111111111111100111010, 
22'b1111111111111100000001, 
22'b0000000000000000011000, 
22'b1111111111111110000000, 
22'b0000000000000010100011, 
22'b1111111111111010110001, 
22'b0000000000000101000001, 
22'b0000000000000011111111, 
22'b0000000000000000010110, 
22'b1111111111111111110100, 
22'b1111111111111011100011, 
22'b1111111111111010101101, 
22'b1111111111111100011001, 
22'b1111111111111101101100, 
22'b1111111111111110111100, 
22'b0000000000000001010001, 
22'b0000000000000111100110, 
22'b1111111111111101110101, 
22'b1111111111111000111010, 
22'b0000000000000111010111, 
22'b1111111111111100011010, 
22'b1111111111111111001000, 
22'b0000000000000001000100, 
22'b0000000000000011010111, 
22'b1111111111111011111010, 
22'b1111111111111100010001, 
22'b1111111111111110011001, 
22'b0000000000000011101111, 
22'b1111111111111100111010, 
22'b0000000000000011001010, 
22'b0000000000000011101011, 
22'b1111111111111010011001, 
22'b0000000000000000001111, 
22'b0000000000000000000111, 
22'b1111111111111110011001, 
22'b1111111111111101100101, 
22'b0000000000000000101100, 
22'b1111111111111110011100, 
22'b0000000000000001110011, 
22'b0000000000000001101100, 
22'b1111111111111010100100, 
22'b1111111111111100010011, 
22'b0000000000000000111010, 
22'b0000000000000011110001, 
22'b1111111111111001000011, 
22'b1111111111110111001110, 
22'b1111111111111100111001, 
22'b1111111111111110100111, 
22'b1111111111111110111100, 
22'b1111111111111111011011, 
22'b1111111111111011011011, 
22'b0000000000000010101100, 
22'b0000000000000010111100, 
22'b1111111111111100111010, 
22'b0000000000000011011010, 
22'b1111111111111111100011, 
22'b1111111111111101110100, 
22'b0000000000000101100010, 
22'b1111111111111100001110, 
22'b1111111111111110110111, 
22'b1111111111111100001100, 
22'b0000000000000001100101, 
22'b0000000000000100100010, 
22'b1111111111111111110001, 
22'b0000000000000010110110, 
22'b1111111111110110111000, 
22'b0000000000000000110110, 
22'b1111111111111100101110, 
22'b1111111111111101011000, 
22'b0000000000000100110100, 
22'b1111111111111010001110, 
22'b0000000000000010101000, 
22'b1111111111111101011110, 
22'b0000000000000000001001, 
22'b0000000000000000001000, 
22'b1111111111111001100101, 
22'b1111111111111111100111, 
22'b0000000000000000111100, 
22'b1111111111111011011011, 
22'b0000000000000001000000, 
22'b0000000000000101000001, 
22'b1111111111111100100010, 
22'b0000000000000011110010, 
22'b1111111111111110001111, 
22'b0000000000000110111100, 
22'b1111111111110101111100, 
22'b1111111111110101100010, 
22'b0000000000000011000110, 
22'b1111111111111101001000, 
22'b0000000000000001010101, 
22'b1111111111111011101111, 
22'b1111111111111110101111, 
22'b0000000000000011101101, 
22'b0000000000000001000100, 
22'b1111111111111111110000, 
22'b0000000000000001000000, 
22'b1111111111111100100101, 
22'b0000000000000100010110, 
22'b1111111111111111110110, 
22'b1111111111111100111010, 
22'b0000000000000010100011, 
22'b1111111111111111000100, 
22'b0000000000000000011101, 
22'b0000000000000011111010, 
22'b1111111111111001001110, 
22'b1111111111111100000011, 
22'b1111111111110101111011, 
22'b0000000000000010000000, 
22'b1111111111111001001010, 
22'b0000000000000011000000, 
22'b0000000000000010011111, 
22'b1111111111111111111110, 
22'b1111111111111011111100, 
22'b1111111111111100101111, 
22'b0000000000000011100111, 
22'b1111111111111111010010, 
22'b1111111111110111111001, 
22'b0000000000000110010111, 
22'b1111111111110111000100, 
22'b1111111111111011001101, 
22'b1111111111111111000010, 
22'b0000000000000000000010, 
22'b1111111111111010010011, 
22'b1111111111111101011011, 
22'b1111111111111111111001, 
22'b1111111111111111011011, 
22'b1111111111111110100000, 
22'b1111111111111111101010, 
22'b1111111111111100010110, 
22'b0000000000000111000111, 
22'b1111111111111110001000, 
22'b0000000000000000111000, 
22'b0000000000000000111010, 
22'b1111111111111110110000, 
22'b0000000000000001010011, 
22'b0000000000000000101110, 
22'b1111111111111110011111, 
22'b1111111111111110100110, 
22'b0000000000000001101101, 
22'b0000000000000000110101, 
22'b0000000000000001011001, 
22'b0000000000000010101101, 
22'b1111111111111011010001, 
22'b0000000000000111110010, 
22'b1111111111111101000011, 
22'b0000000000000001000010, 
22'b1111111111111101010000, 
22'b0000000000000010100110, 
22'b1111111111111010011100, 
22'b1111111111111011100111, 
22'b1111111111111000111011, 
22'b1111111111111110101001, 
22'b1111111111110101100101, 
22'b1111111111111111101100, 
22'b1111111111111100011111, 
22'b1111111111111010010000, 
22'b1111111111111011110001, 
22'b1111111111111101111100, 
22'b1111111111111100010000, 
22'b0000000000000101010001, 
22'b1111111111110101111011, 
22'b0000000000001000010001, 
22'b1111111111111110101111, 
22'b1111111111111011110110, 
22'b1111111111111110101010, 
22'b1111111111111001110110, 
22'b0000000000000001001000, 
22'b0000000000000010110000, 
22'b1111111111111010101101, 
22'b0000000000000001011100, 
22'b1111111111111000100100, 
22'b0000000000000100001000, 
22'b1111111111111001111111, 
22'b0000000000000001011111, 
22'b1111111111111101000100, 
22'b1111111111111110000111, 
22'b0000000000000101100100, 
22'b0000000000000100100101, 
22'b1111111111111100110000, 
22'b0000000000000100011111, 
22'b0000000000000001110000, 
22'b0000000000000001001101, 
22'b0000000000000110110101, 
22'b0000000000000011111010, 
22'b1111111111111100100001, 
22'b1111111111111100000011, 
22'b0000000000000101110001, 
22'b0000000000000101010111, 
22'b0000000000000000011101, 
22'b0000000000000011000010, 
22'b0000000000000001011111, 
22'b0000000000000001011011, 
22'b1111111111111110110001, 
22'b0000000000000100111100, 
22'b1111111111111111000010, 
22'b0000000000000000000111, 
22'b0000000000000001111011, 
22'b0000000000001001100101, 
22'b1111111111111010101101, 
22'b1111111111111101110111, 
22'b0000000000000000001110, 
22'b0000000000000100000000, 
22'b0000000000000100111111, 
22'b1111111111111011000111, 
22'b1111111111111010110001, 
22'b0000000000000000101000, 
22'b0000000000000001110010, 
22'b0000000000000000101001, 
22'b0000000000000001000011, 
22'b0000000000000010010001, 
22'b0000000000000001110101, 
22'b0000000000000100001000, 
22'b1111111111111111110011, 
22'b0000000000000000101101, 
22'b0000000000000100100001, 
22'b1111111111111111101100, 
22'b1111111111111110100010, 
22'b0000000000000001000011, 
22'b1111111111111001100110, 
22'b0000000000000000110000, 
22'b0000000000000010110010, 
22'b1111111111111010111011, 
22'b0000000000000111110110, 
22'b1111111111111111100011, 
22'b0000000000000001111101, 
22'b1111111111111111101010, 
22'b1111111111111110110110, 
22'b1111111111111110100100, 
22'b0000000000000011101110, 
22'b0000000000000111111001, 
22'b0000000000000000000000, 
22'b0000000000000011000011, 
22'b0000000000001000000100, 
22'b1111111111111001111000, 
22'b0000000000000011110001, 
22'b0000000000000100000111, 
22'b1111111111111011110111, 
22'b0000000000000000111110, 
22'b0000000000000100111010, 
22'b0000000000000000011111, 
22'b0000000000000011101001, 
22'b1111111111111111011100, 
22'b0000000000000110111000, 
22'b0000000000000010111101, 
22'b1111111111111101000111, 
22'b1111111111111000011100, 
22'b1111111111111011011100, 
22'b0000000000000001100100, 
22'b0000000000000000011101, 
22'b1111111111111111000011, 
22'b0000000000000010001111, 
22'b0000000000000010110100, 
22'b0000000000000010101001, 
22'b1111111111111000110011, 
22'b0000000000000001011111, 
22'b0000000000000011010011, 
22'b1111111111111001101101, 
22'b1111111111111100101111, 
22'b1111111111111110111011, 
22'b0000000000000110010010, 
22'b0000000000000110101011, 
22'b1111111111111111111001, 
22'b0000000000000011101010, 
22'b1111111111111001101011, 
22'b1111111111111101101011, 
22'b1111111111111101111000, 
22'b1111111111111111001011, 
22'b0000000000000000100101, 
22'b1111111111110111100000, 
22'b0000000000000011101100, 
22'b1111111111111110010110, 
22'b1111111111111110010000, 
22'b1111111111111010100000, 
22'b0000000000000000111011, 
22'b1111111111111111101110, 
22'b0000000000001001011110, 
22'b1111111111111000101111, 
22'b0000000000000010000000, 
22'b0000000000000000001110, 
22'b1111111111111100001011, 
22'b1111111111111101100100, 
22'b0000000000000001010010, 
22'b1111111111111010101100, 
22'b1111111111111100111011, 
22'b1111111111111000111100, 
22'b1111111111111110001101, 
22'b0000000000000011011100, 
22'b0000000000000110011001, 
22'b1111111111111011110110, 
22'b1111111111111110011000, 
22'b0000000000000001001100, 
22'b0000000000000101001010, 
22'b1111111111111101111010, 
22'b1111111111111111111001, 
22'b1111111111111111010100, 
22'b0000000000000101100010, 
22'b1111111111110111011101, 
22'b0000000000000101010110, 
22'b1111111111111100100001, 
22'b1111111111110111110010, 
22'b1111111111111011110000, 
22'b0000000000001000010100, 
22'b1111111111111001011100, 
22'b1111111111111110001001, 
22'b1111111111111000000101, 
22'b0000000000000011000111, 
22'b0000000000000111000011, 
22'b0000000000000111011000, 
22'b1111111111111011111001, 
22'b0000000000000000011000, 
22'b1111111111110111100100, 
22'b0000000000000011011010, 
22'b1111111111111100001000, 
22'b0000000000000100101111, 
22'b0000000000000000001011, 
22'b0000000000000010100001, 
22'b1111111111111100000101, 
22'b1111111111111100110110, 
22'b1111111111111011101110, 
22'b0000000000000001100110, 
22'b0000000000000010001101, 
22'b0000000000000110111111, 
22'b0000000000000001000100, 
22'b1111111111111100001010, 
22'b1111111111111110000111, 
22'b1111111111111001001000, 
22'b0000000000000101010100, 
22'b0000000000000011101101, 
22'b1111111111111010001001, 
22'b1111111111111110011101, 
22'b1111111111110111100110, 
22'b0000000000000101010111, 
22'b1111111111111001100101, 
22'b0000000000000110100011, 
22'b1111111111111011111101, 
22'b0000000000000001100010, 
22'b0000000000000000110110, 
22'b0000000000000101000011, 
22'b1111111111111011011111, 
22'b1111111111111010111111, 
22'b0000000000000101101001, 
22'b1111111111111100110111, 
22'b0000000000000000101000, 
22'b1111111111111010101001, 
22'b0000000000000000011000, 
22'b1111111111111101000010, 
22'b0000000000000011101011, 
22'b1111111111111101101011, 
22'b1111111111111100110101, 
22'b1111111111111101000010, 
22'b0000000000000011001000, 
22'b1111111111111101100100, 
22'b1111111111111110101010, 
22'b0000000000000010100010, 
22'b0000000000000100110111, 
22'b1111111111111000010111, 
22'b0000000000000000100101, 
22'b0000000000000000110111, 
22'b1111111111110111110011, 
22'b1111111111111110110010, 
22'b0000000000000110001010, 
22'b0000000000000011101001, 
22'b1111111111111000111011, 
22'b0000000000000011110110, 
22'b1111111111110010001001, 
22'b1111111111111001011110, 
22'b1111111111111010010101, 
22'b0000000000000000100000, 
22'b1111111111110111010101, 
22'b1111111111111101110011, 
22'b0000000000000000100101, 
22'b1111111111111101000000, 
22'b0000000000000111111110, 
22'b0000000000000001000001, 
22'b0000000000000000010100, 
22'b0000000000000000000000, 
22'b0000000000001001011001, 
22'b1111111111111010011101, 
22'b1111111111111010111111, 
22'b0000000000000001011100, 
22'b0000000000000101010001, 
22'b0000000000000100000011, 
22'b0000000000000100000110, 
22'b1111111111111100010100, 
22'b1111111111111010111100, 
22'b0000000000000000111100, 
22'b1111111111111011101010, 
22'b0000000000000001010111, 
22'b0000000000000001111101, 
22'b0000000000000000101001, 
22'b1111111111111000101110, 
22'b1111111111111000101011, 
22'b1111111111111111001000, 
22'b1111111111111110001111, 
22'b1111111111111110110110, 
22'b1111111111111000001010, 
22'b0000000000000001010111, 
22'b1111111111111101010010, 
22'b1111111111110110101011, 
22'b1111111111111011110101, 
22'b0000000000000101011101, 
22'b1111111111111001111010, 
22'b0000000000000100100111, 
22'b0000000000001000000100, 
22'b0000000000000111111000, 
22'b1111111111111111110000, 
22'b1111111111111010101111, 
22'b0000000000000011011111, 
22'b1111111111111010110001, 
22'b1111111111111101110000, 
22'b0000000000000011001110, 
22'b1111111111111111001000, 
22'b1111111111111110111110, 
22'b1111111111111110110111, 
22'b0000000000000100000111
};
localparam logic signed [21:0] dlBiases [9:0] = {
22'b0000000000000101010100, 
22'b1111111111111111111101, 
22'b1111111111111111111101, 
22'b1111111111111110001000, 
22'b1111111111111110000011, 
22'b1111111111111111010111, 
22'b1111111111111111010011, 
22'b0000000000000010011100, 
22'b1111111111111010001111, 
22'b1111111111111111010111
};
localparam logic signed [21:0] convWeights [0:17] = {
22'b0000000000000011100101, 
22'b0000000000001111011001, 
22'b1111111111111000010111, 
22'b0000000000000010111111, 
22'b0000000000000000011101, 
22'b0000000000010000011011, 
22'b0000000000001100111110, 
22'b0000000000000110011000, 
22'b1111111111111000101100, 
22'b0000000000001011001000, 
22'b1111111111111101001111, 
22'b0000000000000110101110, 
22'b0000000000001111111011, 
22'b0000000000000101000111, 
22'b0000000000001100010000, 
22'b1111111111111111101001, 
22'b0000000000000101110101, 
22'b0000000000000011101001
};
localparam logic signed [21:0] convBiases [1:0] = {
22'b0000000000000000000000, 
22'b0000000000000000000000
};
endpackage