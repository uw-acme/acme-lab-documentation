package data18_7;

localparam logic signed [17:0] dlWeights [0:1279] = {
18'b000000001000001110, 
18'b000000000000010100, 
18'b111111111001110000, 
18'b000000000000001101, 
18'b111111111101111010, 
18'b000000000100010010, 
18'b000000000010000001, 
18'b111111111001101000, 
18'b000000000001011101, 
18'b000000000101010111, 
18'b000000000101011000, 
18'b111111110111101111, 
18'b111111110011110111, 
18'b111111111010100110, 
18'b000000000011000100, 
18'b111111111100001001, 
18'b111111111101100110, 
18'b111111111111000010, 
18'b111111111110011000, 
18'b111111111111111001, 
18'b000000000011110110, 
18'b111111111000010110, 
18'b000000000001101110, 
18'b000000000010100100, 
18'b111111111110111101, 
18'b000000000000001010, 
18'b111111111101111001, 
18'b000000000001000111, 
18'b000000000010000101, 
18'b000000001000000110, 
18'b000000010010010110, 
18'b111111110010010101, 
18'b111111111000001100, 
18'b111111110110101000, 
18'b111111111000100011, 
18'b000000000011111001, 
18'b111111111111001010, 
18'b000000000101001101, 
18'b111111111101101111, 
18'b000000000110100100, 
18'b000000000100111111, 
18'b111111111011101011, 
18'b111111111111011101, 
18'b111111111010100101, 
18'b000000000000001011, 
18'b111111111100111101, 
18'b000000000101100101, 
18'b111111111011001101, 
18'b111111111100011011, 
18'b000000000000010100, 
18'b000000001011101011, 
18'b111111111011011010, 
18'b111111110111110001, 
18'b111111110101010011, 
18'b111111111010110100, 
18'b000000000011000110, 
18'b111111111111010010, 
18'b000000000100000100, 
18'b000000000010000011, 
18'b000000000011010010, 
18'b000000000111110001, 
18'b111111111001101010, 
18'b000000000010000110, 
18'b000000000010001001, 
18'b111111111010100101, 
18'b000000000111010010, 
18'b000000000110110100, 
18'b000000000000000101, 
18'b000000000101100110, 
18'b111111111101011100, 
18'b000000000000000111, 
18'b000000000110101101, 
18'b111111111000111111, 
18'b111111111011000111, 
18'b111111111010111010, 
18'b000000000011001011, 
18'b111111111110101110, 
18'b000000000101101000, 
18'b111111111000100010, 
18'b111111111010001111, 
18'b111111111101100101, 
18'b111111111100101001, 
18'b111111111000110001, 
18'b000000000011010111, 
18'b111111111011101100, 
18'b000000000100010001, 
18'b000000000000000000, 
18'b111111111010100111, 
18'b111111111110001111, 
18'b111111111100011101, 
18'b000000000001001000, 
18'b000000000000100010, 
18'b111111111100100110, 
18'b000000000000111000, 
18'b111111110111000001, 
18'b111111111110010110, 
18'b111111111000010110, 
18'b000000001010000010, 
18'b111111110111101101, 
18'b111111110110010100, 
18'b000000000000101010, 
18'b000000001001100001, 
18'b000000000000001010, 
18'b000000000001000110, 
18'b111111111011001101, 
18'b111111111111001110, 
18'b111111111010010011, 
18'b111111111010101001, 
18'b000000000011011110, 
18'b111111111001110000, 
18'b000000000000111001, 
18'b000000000101010100, 
18'b000000000001000111, 
18'b000000000100000101, 
18'b111111111000000100, 
18'b111111111100110011, 
18'b111111110111100100, 
18'b000000000011100011, 
18'b111111111010101111, 
18'b000000000010000011, 
18'b111111111010000011, 
18'b111111111110001110, 
18'b000000000000100011, 
18'b000000000010011010, 
18'b111111111000011101, 
18'b111111111101111010, 
18'b111111111000100100, 
18'b111111111100110001, 
18'b000000000000000100, 
18'b000000000010101001, 
18'b111111111010110101, 
18'b111111111101111101, 
18'b111111111100101010, 
18'b000000001000111101, 
18'b111111111010011010, 
18'b111111110101110001, 
18'b111111111011010010, 
18'b000000001010001001, 
18'b111111111110010011, 
18'b000000000001100000, 
18'b111111111111100110, 
18'b111111111101011110, 
18'b000000000000011111, 
18'b000000000001100000, 
18'b000000000110011111, 
18'b111111111110101100, 
18'b111111110111100100, 
18'b000000000110100111, 
18'b111111111110010000, 
18'b000000000010001100, 
18'b000000000000101001, 
18'b000000000010101011, 
18'b000000000100101010, 
18'b111111111111101011, 
18'b000000000010100111, 
18'b111111111011010101, 
18'b111111100111111110, 
18'b000000000110011001, 
18'b111111111110100100, 
18'b000000000011001100, 
18'b000000000101000110, 
18'b111111111110001000, 
18'b111111110111101111, 
18'b000000000101111011, 
18'b000000000110111001, 
18'b111111111100100110, 
18'b000000001000000101, 
18'b111111111110001011, 
18'b000000000001010111, 
18'b111111111111011001, 
18'b000000000100101110, 
18'b111111111111100000, 
18'b111111111110001001, 
18'b111111110101000101, 
18'b000000000000100110, 
18'b000000000001110011, 
18'b111111111101010111, 
18'b111111111111001000, 
18'b111111111100011010, 
18'b000000000100101100, 
18'b000000000111100001, 
18'b111111111000100001, 
18'b111111111111011100, 
18'b111111111101000101, 
18'b000000000111100101, 
18'b111111111111101101, 
18'b000000000100011100, 
18'b111111111100011111, 
18'b000000000110010111, 
18'b000000000000001111, 
18'b000000000111100001, 
18'b111111110100111000, 
18'b111111111011010110, 
18'b111111110111100011, 
18'b111111111111110010, 
18'b000000000010111011, 
18'b000000000001010110, 
18'b000000000011010100, 
18'b000000000100111111, 
18'b111111111110100100, 
18'b000000000110100011, 
18'b111111110111101000, 
18'b111111111100100100, 
18'b111111111011101001, 
18'b111111111111111100, 
18'b000000000000010110, 
18'b000000000000000111, 
18'b111111111110111110, 
18'b000000000000101011, 
18'b111111111100110000, 
18'b111111111110001011, 
18'b111111111110101010, 
18'b111111111110100101, 
18'b111111111001011001, 
18'b111111111111100001, 
18'b000000000000110101, 
18'b000000000110101000, 
18'b111111111101000100, 
18'b000000000000011111, 
18'b000000000001011011, 
18'b111111111011101111, 
18'b111111111110011001, 
18'b111111111001110110, 
18'b000000000101111100, 
18'b111111111001101110, 
18'b000000000111101011, 
18'b111111111010010011, 
18'b000000000000100111, 
18'b111111111101010110, 
18'b111111110111011110, 
18'b000000000101000100, 
18'b000000000111010110, 
18'b111111111001111111, 
18'b000000000010001111, 
18'b111111111111010000, 
18'b000000000000011101, 
18'b111111111100101001, 
18'b000000000101000100, 
18'b000000000001111110, 
18'b000000000001100111, 
18'b000000000000000110, 
18'b111111111100101001, 
18'b000000000010101001, 
18'b000000000011110111, 
18'b000000000010100001, 
18'b111111111101011001, 
18'b111111111010101100, 
18'b111111111101111101, 
18'b000000000011110010, 
18'b111111111011010010, 
18'b000000000010011001, 
18'b000000000010001101, 
18'b111111111101100111, 
18'b111111111011111111, 
18'b111111110111101000, 
18'b111111111100101100, 
18'b000000000000010101, 
18'b000000000000000010, 
18'b111111110110010101, 
18'b111111111001011110, 
18'b111111111000000000, 
18'b000000000001011000, 
18'b000000000000111111, 
18'b000000000010110101, 
18'b111111110101010110, 
18'b000000000000101110, 
18'b000000000011100011, 
18'b111111111001011100, 
18'b000000000000010011, 
18'b111111111111001110, 
18'b000000000000111100, 
18'b000000000101111000, 
18'b000000000001101000, 
18'b000000000000111011, 
18'b111111111110111000, 
18'b111111111001100010, 
18'b111111111000111000, 
18'b000000001000011110, 
18'b111111110111001011, 
18'b000000000000101010, 
18'b111111111111101000, 
18'b000000000000010000, 
18'b000000000010110101, 
18'b111111111110010100, 
18'b000000000001000110, 
18'b111111111100100001, 
18'b000000000011010000, 
18'b111111111111111101, 
18'b000000000100100011, 
18'b000000000010111011, 
18'b111111111100100010, 
18'b000000000011101101, 
18'b000000000011101110, 
18'b000000000000001011, 
18'b000000000010110100, 
18'b111111111100111101, 
18'b111111110110010000, 
18'b111111111111011011, 
18'b111111111010100010, 
18'b111111111101110101, 
18'b000000000001001101, 
18'b000000000110011001, 
18'b000000000001100001, 
18'b000000000010111100, 
18'b111111111101110000, 
18'b000000000001010000, 
18'b000000000010101011, 
18'b111111111101111000, 
18'b000000000011001100, 
18'b000000000110011100, 
18'b000000000011111111, 
18'b000000000010011000, 
18'b111111111110110011, 
18'b000000000001100000, 
18'b000000000100101110, 
18'b000000000010101001, 
18'b111111111000011010, 
18'b000000000000100101, 
18'b111111111110101000, 
18'b111111111111110110, 
18'b000000000100001011, 
18'b111111110111011011, 
18'b111111111011100110, 
18'b000000000011011000, 
18'b000000000110111000, 
18'b000000000000100110, 
18'b000000000110111111, 
18'b111111110111110010, 
18'b000000000000010000, 
18'b000000000011110101, 
18'b000000001000111011, 
18'b111111110111100010, 
18'b111111111101010000, 
18'b111111110101110110, 
18'b111111111110000001, 
18'b000000000011001111, 
18'b111111111011111110, 
18'b000000000001011000, 
18'b111111111101001110, 
18'b111111111011010000, 
18'b000000000011110001, 
18'b111111111101010000, 
18'b111111111110011100, 
18'b111111111010000010, 
18'b000000000001001111, 
18'b111111111101110010, 
18'b000000000001111010, 
18'b111111111100101100, 
18'b000000000101000110, 
18'b111111111011100111, 
18'b000000000101000111, 
18'b111111111101101010, 
18'b111111110100110101, 
18'b000000000001100110, 
18'b000000000100110101, 
18'b000000000000010110, 
18'b000000000000110110, 
18'b000000000001000010, 
18'b000000000101001010, 
18'b111111111100111000, 
18'b000000000001011111, 
18'b111111111000001111, 
18'b000000000100000010, 
18'b000000000100100010, 
18'b000000000000100111, 
18'b111111111101111000, 
18'b000000000010100111, 
18'b111111111110000101, 
18'b000000000010001010, 
18'b000000000001000111, 
18'b000000000000000010, 
18'b000000000000110000, 
18'b111111111011001110, 
18'b000000000001100000, 
18'b111111111110100111, 
18'b000000000001001111, 
18'b000000000110101001, 
18'b000000000100010110, 
18'b111111111111010010, 
18'b111111111001101010, 
18'b000000000011100100, 
18'b111111111000101010, 
18'b111111111101111111, 
18'b111111111100111101, 
18'b111111111111110111, 
18'b000000000101011110, 
18'b111111111110010110, 
18'b000000000000000101, 
18'b000000000111110000, 
18'b111111111110100010, 
18'b111111111110100010, 
18'b111111111101111001, 
18'b111111111111011000, 
18'b000000000100001001, 
18'b111111111010010000, 
18'b111111111101001111, 
18'b111111111101010101, 
18'b111111111001110101, 
18'b111111111011110001, 
18'b111111110111101001, 
18'b111111111100101101, 
18'b111111111100111001, 
18'b111111110111111110, 
18'b000000000110001100, 
18'b111111111001111111, 
18'b000000000010001100, 
18'b111111111010101111, 
18'b111111111010110010, 
18'b000000000011110111, 
18'b000000000000000111, 
18'b111111111010010100, 
18'b000000000001011101, 
18'b111111111001011100, 
18'b000000000101001001, 
18'b000000000010010001, 
18'b111111111101101000, 
18'b111111111011110111, 
18'b111111111100000110, 
18'b000000000011001110, 
18'b111111111010000000, 
18'b000000000000010101, 
18'b000000000101001001, 
18'b000000000010110000, 
18'b000000000011011010, 
18'b111111111010011001, 
18'b000000000110011110, 
18'b000000000100111011, 
18'b000000000000110010, 
18'b000000000111010000, 
18'b000000000000111010, 
18'b111111110111001111, 
18'b000000000110110000, 
18'b000000000010100111, 
18'b000000000101100110, 
18'b111111111000111000, 
18'b111111111110100111, 
18'b000000000001110011, 
18'b111111111010011101, 
18'b111111111011001001, 
18'b111111111011011100, 
18'b111111111100101110, 
18'b000000000111010100, 
18'b000000000000011011, 
18'b000000000011010001, 
18'b000000000000011001, 
18'b000000000110000101, 
18'b000000000101110001, 
18'b111111111000011111, 
18'b111111111010110000, 
18'b000000000100011010, 
18'b111111111011110111, 
18'b111111111110110000, 
18'b111111111110110001, 
18'b000000000100000111, 
18'b000000000001100011, 
18'b111111111111101110, 
18'b111111111010101011, 
18'b000000000100111101, 
18'b111111111110010101, 
18'b000000000101011100, 
18'b000000000001111010, 
18'b000000000010101010, 
18'b111111111101111100, 
18'b000000000000100011, 
18'b000000000101011100, 
18'b111111111110111011, 
18'b111111111111101000, 
18'b111111111111010001, 
18'b111111111011001111, 
18'b000000001000000010, 
18'b000000000001001101, 
18'b111111111100001011, 
18'b111111111111010101, 
18'b000000000001110001, 
18'b111111111110100111, 
18'b111111111110100010, 
18'b000000000001001000, 
18'b000000000110010110, 
18'b000000000011100011, 
18'b000000000101101100, 
18'b000000000001111110, 
18'b111111111011010000, 
18'b000000000001010000, 
18'b111111111011010001, 
18'b111111111101010100, 
18'b111111111100001001, 
18'b000000000000000010, 
18'b000000000000101100, 
18'b000000000010101110, 
18'b000000000001100111, 
18'b000000000010000010, 
18'b111111110110011100, 
18'b111111111011000000, 
18'b111111111111000011, 
18'b000000000000111000, 
18'b000000000111101101, 
18'b000000000111100011, 
18'b111111110111100110, 
18'b111111111110111111, 
18'b000000000100001001, 
18'b000000000110101100, 
18'b111111110111100110, 
18'b111111111011010010, 
18'b000000000000111000, 
18'b000000000100101101, 
18'b111111111101000110, 
18'b111111111101110110, 
18'b111111111110010011, 
18'b111111111111101011, 
18'b000000000110101101, 
18'b000000000101010011, 
18'b111111111111011011, 
18'b111111111101101100, 
18'b000000000100101100, 
18'b000000000010010001, 
18'b000000000100010101, 
18'b111111111111001111, 
18'b111111111100001111, 
18'b111111111110001100, 
18'b111111111111001000, 
18'b111111111001010000, 
18'b000000000001011011, 
18'b111111111001100001, 
18'b000000000011001111, 
18'b111111111111000011, 
18'b111111111111001010, 
18'b000000000100000110, 
18'b000000000000100111, 
18'b111111111111010110, 
18'b000000000010101101, 
18'b000000000010000110, 
18'b000000000001101111, 
18'b000000000000110111, 
18'b000000000011000000, 
18'b111111111011111010, 
18'b000000001000000101, 
18'b000000000011111101, 
18'b111111110111010011, 
18'b000000000000100101, 
18'b111111111001000011, 
18'b111111111000110000, 
18'b111111110110101111, 
18'b111111111110010100, 
18'b111111111101010110, 
18'b111111111100000111, 
18'b000000000010110110, 
18'b000000000000100000, 
18'b111111111001111101, 
18'b000000000001010010, 
18'b111111111100001101, 
18'b111111111100100001, 
18'b111111111101000000, 
18'b111111111101111011, 
18'b111111111100110001, 
18'b000000000000100010, 
18'b111111111110010011, 
18'b000000000100101100, 
18'b111111111100000010, 
18'b000000000001101100, 
18'b000000000000110011, 
18'b000000000010110010, 
18'b000000000110110011, 
18'b000000000000000011, 
18'b111111111011101010, 
18'b111111111101000001, 
18'b000000000011100101, 
18'b000000000100011101, 
18'b111111110101111010, 
18'b000000000010011011, 
18'b000000000000100111, 
18'b111111110111010100, 
18'b000000000101101011, 
18'b111111111101100010, 
18'b000000000000001001, 
18'b111111111011011100, 
18'b000000000101100001, 
18'b000000000011111001, 
18'b111111110100110101, 
18'b000000000100011100, 
18'b000000000010111111, 
18'b000000000010110010, 
18'b000000001001010011, 
18'b000000000010100111, 
18'b000000000101000101, 
18'b111111111011000110, 
18'b000000000001001001, 
18'b111111111110001001, 
18'b000000000010001001, 
18'b000000000111011000, 
18'b000000000011101101, 
18'b111111110101110100, 
18'b000000000101001101, 
18'b111111111101101100, 
18'b000000000001011011, 
18'b111111111011111010, 
18'b111111111010010010, 
18'b000000000001000110, 
18'b000000000011110001, 
18'b000000000001111011, 
18'b111111111110001100, 
18'b111111110110110001, 
18'b000000000010010100, 
18'b000000000000110111, 
18'b000000000100101000, 
18'b000000000000001100, 
18'b000000000001000101, 
18'b000000000100111010, 
18'b000000000100010001, 
18'b111111111101101101, 
18'b000000000011011100, 
18'b111111111011111011, 
18'b111111111011111101, 
18'b111111111101010001, 
18'b000000000101100100, 
18'b111111111100001110, 
18'b111111111010011111, 
18'b000000000000111011, 
18'b000000000011011110, 
18'b000000000100010010, 
18'b111111111100111010, 
18'b111111110111011100, 
18'b111111110111001110, 
18'b000000000011110100, 
18'b000000000000011111, 
18'b000000000101011100, 
18'b000000000100011011, 
18'b000000000011101110, 
18'b000000000101110000, 
18'b111111111101001110, 
18'b111111111111100000, 
18'b000000000001011011, 
18'b000000000010010101, 
18'b000000000100111001, 
18'b000000000101011100, 
18'b000000000110100001, 
18'b111111111011110011, 
18'b000000000000000010, 
18'b000000000110101001, 
18'b000000000100110111, 
18'b000000000100100010, 
18'b111111111111100111, 
18'b111111111010111111, 
18'b111111111110101000, 
18'b111111111110110100, 
18'b111111111011110001, 
18'b111111111000001000, 
18'b000000000100001111, 
18'b000000000011110000, 
18'b000000000101000011, 
18'b000000000000000100, 
18'b111111111100111101, 
18'b111111111110101110, 
18'b111111111100001101, 
18'b000000000000111101, 
18'b000000000000000101, 
18'b000000000101111010, 
18'b000000000010100110, 
18'b111111110111000101, 
18'b111111111011011100, 
18'b111111111010010110, 
18'b111111111111110010, 
18'b111111111000110000, 
18'b111111111110011110, 
18'b111111111101101000, 
18'b000000000001101111, 
18'b000000000000010011, 
18'b000000000001000111, 
18'b111111110110011011, 
18'b111111111111101000, 
18'b000000000100010100, 
18'b000000000110110001, 
18'b111111111111010101, 
18'b111111111000011111, 
18'b000000000011110011, 
18'b111111111110001100, 
18'b000000000101101010, 
18'b111111111111110100, 
18'b111111110110111111, 
18'b111111111101000011, 
18'b000000000000101100, 
18'b111111111000100111, 
18'b111111111111010101, 
18'b000000000101101001, 
18'b111111111101101000, 
18'b111111111111101011, 
18'b000000000101011111, 
18'b000000000001110110, 
18'b111111111101101110, 
18'b000000000101110001, 
18'b111111111101110001, 
18'b000000000010011001, 
18'b000000000000011011, 
18'b111111111001110100, 
18'b000000000101000010, 
18'b111111111100110110, 
18'b000000000000010011, 
18'b000000000000101001, 
18'b111111111101001111, 
18'b111111111110011001, 
18'b000000000011100010, 
18'b000000000000000100, 
18'b000000000001011010, 
18'b000000000010011010, 
18'b111111111100011101, 
18'b000000000001110101, 
18'b111111111010101101, 
18'b111111111111110111, 
18'b111111111100110110, 
18'b111111111100101000, 
18'b111111111011001001, 
18'b000000000000110000, 
18'b000000000010101000, 
18'b000000000001011110, 
18'b111111111101100001, 
18'b111111111011010100, 
18'b000000000101010011, 
18'b111111111100111110, 
18'b000000000000000010, 
18'b000000000110011110, 
18'b000000000000001000, 
18'b111111111001100101, 
18'b000000000100011010, 
18'b111111111011100110, 
18'b000000000010111011, 
18'b000000000001111110, 
18'b000000000010000010, 
18'b000000000100001110, 
18'b111111111011000011, 
18'b000000000001100101, 
18'b111111111100110001, 
18'b111111111010001011, 
18'b000000000011011100, 
18'b111111111001110101, 
18'b000000000101101011, 
18'b000000000001000101, 
18'b111111111101110000, 
18'b111111111001100100, 
18'b111111111101001111, 
18'b000000000101010011, 
18'b111111111100000110, 
18'b000000000000010100, 
18'b111111111101010010, 
18'b000000000110000001, 
18'b111111111110111100, 
18'b000000000000100110, 
18'b000000000011000010, 
18'b111111111100110101, 
18'b111111111100011000, 
18'b000000000001100000, 
18'b000000000000110011, 
18'b111111111000101000, 
18'b000000000110110100, 
18'b111111111110100101, 
18'b000000000110010100, 
18'b000000000011100010, 
18'b000000000011001001, 
18'b111111111011100001, 
18'b111111111110100001, 
18'b111111111110100000, 
18'b111111111101110000, 
18'b111111111111010110, 
18'b000000000011100010, 
18'b111111111100000111, 
18'b000000000011001100, 
18'b000000000000101110, 
18'b000000000001000101, 
18'b000000000011010011, 
18'b000000000101000010, 
18'b000000000010101010, 
18'b111111111100010000, 
18'b000000000001110101, 
18'b111111111000011111, 
18'b000000000010001001, 
18'b111111111101101000, 
18'b000000000011000101, 
18'b111111111101001001, 
18'b111111111100100111, 
18'b000000000010101010, 
18'b111111111011000110, 
18'b111111111100111111, 
18'b111111111010100110, 
18'b000000000000111011, 
18'b111111111100011010, 
18'b000000000111001101, 
18'b111111111111010011, 
18'b111111111100010001, 
18'b111111111111111000, 
18'b000000000010100100, 
18'b000000000010100001, 
18'b000000000101011111, 
18'b111111111101011111, 
18'b111111111010000000, 
18'b000000000000011010, 
18'b111111111011110110, 
18'b111111111101011100, 
18'b111111111001000000, 
18'b000000000011011000, 
18'b000000001000011010, 
18'b000000000011001110, 
18'b000000000101001110, 
18'b111111111111110010, 
18'b111111111100011001, 
18'b000000000100100000, 
18'b111111111110000111, 
18'b000000000101000110, 
18'b111111111101100110, 
18'b000000000001011101, 
18'b111111111010001100, 
18'b000000001000110001, 
18'b000000000111100100, 
18'b111111111100100111, 
18'b111111110101110011, 
18'b000000000000101110, 
18'b111111111011000110, 
18'b000000001000000111, 
18'b111111111111000001, 
18'b111111111100110110, 
18'b000000000000110101, 
18'b111111111100011000, 
18'b111111111100101011, 
18'b111111111101110110, 
18'b111111110110011111, 
18'b000000000000111100, 
18'b111111110110101001, 
18'b111111111101010101, 
18'b000000000000110110, 
18'b000000000010111010, 
18'b111111111100011110, 
18'b111111111111011100, 
18'b000000000001010000, 
18'b111111111101101101, 
18'b111111110101010001, 
18'b111111111101101011, 
18'b000000000001101010, 
18'b000000000001001011, 
18'b000000000010010101, 
18'b000000000010100010, 
18'b111111110111011100, 
18'b111111111101000001, 
18'b000000000101100011, 
18'b111111111001110011, 
18'b111111111101110001, 
18'b000000000111011101, 
18'b111111111100110001, 
18'b000000000000001101, 
18'b111111111100111001, 
18'b000000000001000010, 
18'b111111111110101111, 
18'b111111111101110011, 
18'b000000000101111100, 
18'b111111111001111110, 
18'b111111111101110011, 
18'b000000000100100101, 
18'b000000000101110100, 
18'b111111111110010101, 
18'b000000000010000101, 
18'b111111111110110000, 
18'b111111110111010001, 
18'b111111111101111000, 
18'b000000000001001001, 
18'b111111111100111000, 
18'b111111111111110000, 
18'b111111111110000000, 
18'b111111111100111001, 
18'b000000000100110101, 
18'b111111111100111010, 
18'b111111111100000001, 
18'b000000000000011000, 
18'b111111111110000000, 
18'b000000000010100011, 
18'b111111111010110001, 
18'b000000000101000001, 
18'b000000000011111111, 
18'b000000000000010110, 
18'b111111111111110100, 
18'b111111111011100011, 
18'b111111111010101101, 
18'b111111111100011001, 
18'b111111111101101100, 
18'b111111111110111100, 
18'b000000000001010001, 
18'b000000000111100110, 
18'b111111111101110101, 
18'b111111111000111010, 
18'b000000000111010111, 
18'b111111111100011010, 
18'b111111111111001000, 
18'b000000000001000100, 
18'b000000000011010111, 
18'b111111111011111010, 
18'b111111111100010001, 
18'b111111111110011001, 
18'b000000000011101111, 
18'b111111111100111010, 
18'b000000000011001010, 
18'b000000000011101011, 
18'b111111111010011001, 
18'b000000000000001111, 
18'b000000000000000111, 
18'b111111111110011001, 
18'b111111111101100101, 
18'b000000000000101100, 
18'b111111111110011100, 
18'b000000000001110011, 
18'b000000000001101100, 
18'b111111111010100100, 
18'b111111111100010011, 
18'b000000000000111010, 
18'b000000000011110001, 
18'b111111111001000011, 
18'b111111110111001110, 
18'b111111111100111001, 
18'b111111111110100111, 
18'b111111111110111100, 
18'b111111111111011011, 
18'b111111111011011011, 
18'b000000000010101100, 
18'b000000000010111100, 
18'b111111111100111010, 
18'b000000000011011010, 
18'b111111111111100011, 
18'b111111111101110100, 
18'b000000000101100010, 
18'b111111111100001110, 
18'b111111111110110111, 
18'b111111111100001100, 
18'b000000000001100101, 
18'b000000000100100010, 
18'b111111111111110001, 
18'b000000000010110110, 
18'b111111110110111000, 
18'b000000000000110110, 
18'b111111111100101110, 
18'b111111111101011000, 
18'b000000000100110100, 
18'b111111111010001110, 
18'b000000000010101000, 
18'b111111111101011110, 
18'b000000000000001001, 
18'b000000000000001000, 
18'b111111111001100101, 
18'b111111111111100111, 
18'b000000000000111100, 
18'b111111111011011011, 
18'b000000000001000000, 
18'b000000000101000001, 
18'b111111111100100010, 
18'b000000000011110010, 
18'b111111111110001111, 
18'b000000000110111100, 
18'b111111110101111100, 
18'b111111110101100010, 
18'b000000000011000110, 
18'b111111111101001000, 
18'b000000000001010101, 
18'b111111111011101111, 
18'b111111111110101111, 
18'b000000000011101101, 
18'b000000000001000100, 
18'b111111111111110000, 
18'b000000000001000000, 
18'b111111111100100101, 
18'b000000000100010110, 
18'b111111111111110110, 
18'b111111111100111010, 
18'b000000000010100011, 
18'b111111111111000100, 
18'b000000000000011101, 
18'b000000000011111010, 
18'b111111111001001110, 
18'b111111111100000011, 
18'b111111110101111011, 
18'b000000000010000000, 
18'b111111111001001010, 
18'b000000000011000000, 
18'b000000000010011111, 
18'b111111111111111110, 
18'b111111111011111100, 
18'b111111111100101111, 
18'b000000000011100111, 
18'b111111111111010010, 
18'b111111110111111001, 
18'b000000000110010111, 
18'b111111110111000100, 
18'b111111111011001101, 
18'b111111111111000010, 
18'b000000000000000010, 
18'b111111111010010011, 
18'b111111111101011011, 
18'b111111111111111001, 
18'b111111111111011011, 
18'b111111111110100000, 
18'b111111111111101010, 
18'b111111111100010110, 
18'b000000000111000111, 
18'b111111111110001000, 
18'b000000000000111000, 
18'b000000000000111010, 
18'b111111111110110000, 
18'b000000000001010011, 
18'b000000000000101110, 
18'b111111111110011111, 
18'b111111111110100110, 
18'b000000000001101101, 
18'b000000000000110101, 
18'b000000000001011001, 
18'b000000000010101101, 
18'b111111111011010001, 
18'b000000000111110010, 
18'b111111111101000011, 
18'b000000000001000010, 
18'b111111111101010000, 
18'b000000000010100110, 
18'b111111111010011100, 
18'b111111111011100111, 
18'b111111111000111011, 
18'b111111111110101001, 
18'b111111110101100101, 
18'b111111111111101100, 
18'b111111111100011111, 
18'b111111111010010000, 
18'b111111111011110001, 
18'b111111111101111100, 
18'b111111111100010000, 
18'b000000000101010001, 
18'b111111110101111011, 
18'b000000001000010001, 
18'b111111111110101111, 
18'b111111111011110110, 
18'b111111111110101010, 
18'b111111111001110110, 
18'b000000000001001000, 
18'b000000000010110000, 
18'b111111111010101101, 
18'b000000000001011100, 
18'b111111111000100100, 
18'b000000000100001000, 
18'b111111111001111111, 
18'b000000000001011111, 
18'b111111111101000100, 
18'b111111111110000111, 
18'b000000000101100100, 
18'b000000000100100101, 
18'b111111111100110000, 
18'b000000000100011111, 
18'b000000000001110000, 
18'b000000000001001101, 
18'b000000000110110101, 
18'b000000000011111010, 
18'b111111111100100001, 
18'b111111111100000011, 
18'b000000000101110001, 
18'b000000000101010111, 
18'b000000000000011101, 
18'b000000000011000010, 
18'b000000000001011111, 
18'b000000000001011011, 
18'b111111111110110001, 
18'b000000000100111100, 
18'b111111111111000010, 
18'b000000000000000111, 
18'b000000000001111011, 
18'b000000001001100101, 
18'b111111111010101101, 
18'b111111111101110111, 
18'b000000000000001110, 
18'b000000000100000000, 
18'b000000000100111111, 
18'b111111111011000111, 
18'b111111111010110001, 
18'b000000000000101000, 
18'b000000000001110010, 
18'b000000000000101001, 
18'b000000000001000011, 
18'b000000000010010001, 
18'b000000000001110101, 
18'b000000000100001000, 
18'b111111111111110011, 
18'b000000000000101101, 
18'b000000000100100001, 
18'b111111111111101100, 
18'b111111111110100010, 
18'b000000000001000011, 
18'b111111111001100110, 
18'b000000000000110000, 
18'b000000000010110010, 
18'b111111111010111011, 
18'b000000000111110110, 
18'b111111111111100011, 
18'b000000000001111101, 
18'b111111111111101010, 
18'b111111111110110110, 
18'b111111111110100100, 
18'b000000000011101110, 
18'b000000000111111001, 
18'b000000000000000000, 
18'b000000000011000011, 
18'b000000001000000100, 
18'b111111111001111000, 
18'b000000000011110001, 
18'b000000000100000111, 
18'b111111111011110111, 
18'b000000000000111110, 
18'b000000000100111010, 
18'b000000000000011111, 
18'b000000000011101001, 
18'b111111111111011100, 
18'b000000000110111000, 
18'b000000000010111101, 
18'b111111111101000111, 
18'b111111111000011100, 
18'b111111111011011100, 
18'b000000000001100100, 
18'b000000000000011101, 
18'b111111111111000011, 
18'b000000000010001111, 
18'b000000000010110100, 
18'b000000000010101001, 
18'b111111111000110011, 
18'b000000000001011111, 
18'b000000000011010011, 
18'b111111111001101101, 
18'b111111111100101111, 
18'b111111111110111011, 
18'b000000000110010010, 
18'b000000000110101011, 
18'b111111111111111001, 
18'b000000000011101010, 
18'b111111111001101011, 
18'b111111111101101011, 
18'b111111111101111000, 
18'b111111111111001011, 
18'b000000000000100101, 
18'b111111110111100000, 
18'b000000000011101100, 
18'b111111111110010110, 
18'b111111111110010000, 
18'b111111111010100000, 
18'b000000000000111011, 
18'b111111111111101110, 
18'b000000001001011110, 
18'b111111111000101111, 
18'b000000000010000000, 
18'b000000000000001110, 
18'b111111111100001011, 
18'b111111111101100100, 
18'b000000000001010010, 
18'b111111111010101100, 
18'b111111111100111011, 
18'b111111111000111100, 
18'b111111111110001101, 
18'b000000000011011100, 
18'b000000000110011001, 
18'b111111111011110110, 
18'b111111111110011000, 
18'b000000000001001100, 
18'b000000000101001010, 
18'b111111111101111010, 
18'b111111111111111001, 
18'b111111111111010100, 
18'b000000000101100010, 
18'b111111110111011101, 
18'b000000000101010110, 
18'b111111111100100001, 
18'b111111110111110010, 
18'b111111111011110000, 
18'b000000001000010100, 
18'b111111111001011100, 
18'b111111111110001001, 
18'b111111111000000101, 
18'b000000000011000111, 
18'b000000000111000011, 
18'b000000000111011000, 
18'b111111111011111001, 
18'b000000000000011000, 
18'b111111110111100100, 
18'b000000000011011010, 
18'b111111111100001000, 
18'b000000000100101111, 
18'b000000000000001011, 
18'b000000000010100001, 
18'b111111111100000101, 
18'b111111111100110110, 
18'b111111111011101110, 
18'b000000000001100110, 
18'b000000000010001101, 
18'b000000000110111111, 
18'b000000000001000100, 
18'b111111111100001010, 
18'b111111111110000111, 
18'b111111111001001000, 
18'b000000000101010100, 
18'b000000000011101101, 
18'b111111111010001001, 
18'b111111111110011101, 
18'b111111110111100110, 
18'b000000000101010111, 
18'b111111111001100101, 
18'b000000000110100011, 
18'b111111111011111101, 
18'b000000000001100010, 
18'b000000000000110110, 
18'b000000000101000011, 
18'b111111111011011111, 
18'b111111111010111111, 
18'b000000000101101001, 
18'b111111111100110111, 
18'b000000000000101000, 
18'b111111111010101001, 
18'b000000000000011000, 
18'b111111111101000010, 
18'b000000000011101011, 
18'b111111111101101011, 
18'b111111111100110101, 
18'b111111111101000010, 
18'b000000000011001000, 
18'b111111111101100100, 
18'b111111111110101010, 
18'b000000000010100010, 
18'b000000000100110111, 
18'b111111111000010111, 
18'b000000000000100101, 
18'b000000000000110111, 
18'b111111110111110011, 
18'b111111111110110010, 
18'b000000000110001010, 
18'b000000000011101001, 
18'b111111111000111011, 
18'b000000000011110110, 
18'b111111110010001001, 
18'b111111111001011110, 
18'b111111111010010101, 
18'b000000000000100000, 
18'b111111110111010101, 
18'b111111111101110011, 
18'b000000000000100101, 
18'b111111111101000000, 
18'b000000000111111110, 
18'b000000000001000001, 
18'b000000000000010100, 
18'b000000000000000000, 
18'b000000001001011001, 
18'b111111111010011101, 
18'b111111111010111111, 
18'b000000000001011100, 
18'b000000000101010001, 
18'b000000000100000011, 
18'b000000000100000110, 
18'b111111111100010100, 
18'b111111111010111100, 
18'b000000000000111100, 
18'b111111111011101010, 
18'b000000000001010111, 
18'b000000000001111101, 
18'b000000000000101001, 
18'b111111111000101110, 
18'b111111111000101011, 
18'b111111111111001000, 
18'b111111111110001111, 
18'b111111111110110110, 
18'b111111111000001010, 
18'b000000000001010111, 
18'b111111111101010010, 
18'b111111110110101011, 
18'b111111111011110101, 
18'b000000000101011101, 
18'b111111111001111010, 
18'b000000000100100111, 
18'b000000001000000100, 
18'b000000000111111000, 
18'b111111111111110000, 
18'b111111111010101111, 
18'b000000000011011111, 
18'b111111111010110001, 
18'b111111111101110000, 
18'b000000000011001110, 
18'b111111111111001000, 
18'b111111111110111110, 
18'b111111111110110111, 
18'b000000000100000111
};

localparam logic signed [17:0] dlBiases [9:0] = {
18'b000000000101010100, 
18'b111111111111111101, 
18'b111111111111111101, 
18'b111111111110001000, 
18'b111111111110000011, 
18'b111111111111010111, 
18'b111111111111010011, 
18'b000000000010011100, 
18'b111111111010001111, 
18'b111111111111010111
};

localparam logic signed [17:0] convWeights [0:17] = {
18'b000000000011100101, 
18'b000000001111011001, 
18'b111111111000010111, 
18'b000000000010111111, 
18'b000000000000011101, 
18'b000000010000011011, 
18'b000000001100111110, 
18'b000000000110011000, 
18'b111111111000101100, 
18'b000000001011001000, 
18'b111111111101001111, 
18'b000000000110101110, 
18'b000000001111111011, 
18'b000000000101000111, 
18'b000000001100010000, 
18'b111111111111101001, 
18'b000000000101110101, 
18'b000000000011101001
};

localparam logic signed [17:0] convBiases [1:0] = {
18'b000000000000000000, 
18'b000000000000000000
};
endpackage




