package data8_6;

localparam logic signed [7:0] dlWeights [0:1279] = {
8'b00010000, 
8'b00000000, 
8'b11110011, 
8'b00000000, 
8'b11111011, 
8'b00001000, 
8'b00000100, 
8'b11110011, 
8'b00000010, 
8'b00001010, 
8'b00001010, 
8'b11101111, 
8'b11100111, 
8'b11110101, 
8'b00000110, 
8'b11111000, 
8'b11111011, 
8'b11111110, 
8'b11111100, 
8'b11111111, 
8'b00000111, 
8'b11110000, 
8'b00000011, 
8'b00000101, 
8'b11111101, 
8'b00000000, 
8'b11111011, 
8'b00000010, 
8'b00000100, 
8'b00010000, 
8'b00100100, 
8'b11100100, 
8'b11110000, 
8'b11101101, 
8'b11110001, 
8'b00000111, 
8'b11111110, 
8'b00001010, 
8'b11111011, 
8'b00001101, 
8'b00001001, 
8'b11110111, 
8'b11111110, 
8'b11110101, 
8'b00000000, 
8'b11111001, 
8'b00001011, 
8'b11110110, 
8'b11111000, 
8'b00000000, 
8'b00010111, 
8'b11110110, 
8'b11101111, 
8'b11101010, 
8'b11110101, 
8'b00000110, 
8'b11111110, 
8'b00001000, 
8'b00000100, 
8'b00000110, 
8'b00001111, 
8'b11110011, 
8'b00000100, 
8'b00000100, 
8'b11110101, 
8'b00001110, 
8'b00001101, 
8'b00000000, 
8'b00001011, 
8'b11111010, 
8'b00000000, 
8'b00001101, 
8'b11110001, 
8'b11110110, 
8'b11110101, 
8'b00000110, 
8'b11111101, 
8'b00001011, 
8'b11110001, 
8'b11110100, 
8'b11111011, 
8'b11111001, 
8'b11110001, 
8'b00000110, 
8'b11110111, 
8'b00001000, 
8'b00000000, 
8'b11110101, 
8'b11111100, 
8'b11111000, 
8'b00000010, 
8'b00000001, 
8'b11111001, 
8'b00000001, 
8'b11101110, 
8'b11111100, 
8'b11110000, 
8'b00010100, 
8'b11101111, 
8'b11101100, 
8'b00000001, 
8'b00010011, 
8'b00000000, 
8'b00000010, 
8'b11110110, 
8'b11111110, 
8'b11110100, 
8'b11110101, 
8'b00000110, 
8'b11110011, 
8'b00000001, 
8'b00001010, 
8'b00000010, 
8'b00001000, 
8'b11110000, 
8'b11111001, 
8'b11101111, 
8'b00000111, 
8'b11110101, 
8'b00000100, 
8'b11110100, 
8'b11111100, 
8'b00000001, 
8'b00000100, 
8'b11110000, 
8'b11111011, 
8'b11110001, 
8'b11111001, 
8'b00000000, 
8'b00000101, 
8'b11110101, 
8'b11111011, 
8'b11111001, 
8'b00010001, 
8'b11110100, 
8'b11101011, 
8'b11110110, 
8'b00010100, 
8'b11111100, 
8'b00000011, 
8'b11111111, 
8'b11111010, 
8'b00000000, 
8'b00000011, 
8'b00001100, 
8'b11111101, 
8'b11101111, 
8'b00001101, 
8'b11111100, 
8'b00000100, 
8'b00000001, 
8'b00000101, 
8'b00001001, 
8'b11111111, 
8'b00000101, 
8'b11110110, 
8'b11001111, 
8'b00001100, 
8'b11111101, 
8'b00000110, 
8'b00001010, 
8'b11111100, 
8'b11101111, 
8'b00001011, 
8'b00001101, 
8'b11111001, 
8'b00010000, 
8'b11111100, 
8'b00000010, 
8'b11111110, 
8'b00001001, 
8'b11111111, 
8'b11111100, 
8'b11101010, 
8'b00000001, 
8'b00000011, 
8'b11111010, 
8'b11111110, 
8'b11111000, 
8'b00001001, 
8'b00001111, 
8'b11110001, 
8'b11111110, 
8'b11111010, 
8'b00001111, 
8'b11111111, 
8'b00001000, 
8'b11111000, 
8'b00001100, 
8'b00000000, 
8'b00001111, 
8'b11101001, 
8'b11110110, 
8'b11101111, 
8'b11111111, 
8'b00000101, 
8'b00000010, 
8'b00000110, 
8'b00001001, 
8'b11111101, 
8'b00001101, 
8'b11101111, 
8'b11111001, 
8'b11110111, 
8'b11111111, 
8'b00000000, 
8'b00000000, 
8'b11111101, 
8'b00000001, 
8'b11111001, 
8'b11111100, 
8'b11111101, 
8'b11111101, 
8'b11110010, 
8'b11111111, 
8'b00000001, 
8'b00001101, 
8'b11111010, 
8'b00000000, 
8'b00000010, 
8'b11110111, 
8'b11111100, 
8'b11110011, 
8'b00001011, 
8'b11110011, 
8'b00001111, 
8'b11110100, 
8'b00000001, 
8'b11111010, 
8'b11101110, 
8'b00001010, 
8'b00001110, 
8'b11110011, 
8'b00000100, 
8'b11111110, 
8'b00000000, 
8'b11111001, 
8'b00001010, 
8'b00000011, 
8'b00000011, 
8'b00000000, 
8'b11111001, 
8'b00000101, 
8'b00000111, 
8'b00000101, 
8'b11111010, 
8'b11110101, 
8'b11111011, 
8'b00000111, 
8'b11110110, 
8'b00000100, 
8'b00000100, 
8'b11111011, 
8'b11110111, 
8'b11101111, 
8'b11111001, 
8'b00000000, 
8'b00000000, 
8'b11101100, 
8'b11110010, 
8'b11110000, 
8'b00000010, 
8'b00000001, 
8'b00000101, 
8'b11101010, 
8'b00000001, 
8'b00000111, 
8'b11110010, 
8'b00000000, 
8'b11111110, 
8'b00000001, 
8'b00001011, 
8'b00000011, 
8'b00000001, 
8'b11111101, 
8'b11110011, 
8'b11110001, 
8'b00010000, 
8'b11101110, 
8'b00000001, 
8'b11111111, 
8'b00000000, 
8'b00000101, 
8'b11111100, 
8'b00000010, 
8'b11111001, 
8'b00000110, 
8'b11111111, 
8'b00001001, 
8'b00000101, 
8'b11111001, 
8'b00000111, 
8'b00000111, 
8'b00000000, 
8'b00000101, 
8'b11111001, 
8'b11101100, 
8'b11111110, 
8'b11110101, 
8'b11111011, 
8'b00000010, 
8'b00001100, 
8'b00000011, 
8'b00000101, 
8'b11111011, 
8'b00000010, 
8'b00000101, 
8'b11111011, 
8'b00000110, 
8'b00001100, 
8'b00000111, 
8'b00000100, 
8'b11111101, 
8'b00000011, 
8'b00001001, 
8'b00000101, 
8'b11110000, 
8'b00000001, 
8'b11111101, 
8'b11111111, 
8'b00001000, 
8'b11101110, 
8'b11110111, 
8'b00000110, 
8'b00001101, 
8'b00000001, 
8'b00001101, 
8'b11101111, 
8'b00000000, 
8'b00000111, 
8'b00010001, 
8'b11101111, 
8'b11111010, 
8'b11101011, 
8'b11111100, 
8'b00000110, 
8'b11110111, 
8'b00000010, 
8'b11111010, 
8'b11110110, 
8'b00000111, 
8'b11111010, 
8'b11111100, 
8'b11110100, 
8'b00000010, 
8'b11111011, 
8'b00000011, 
8'b11111001, 
8'b00001010, 
8'b11110111, 
8'b00001010, 
8'b11111011, 
8'b11101001, 
8'b00000011, 
8'b00001001, 
8'b00000000, 
8'b00000001, 
8'b00000010, 
8'b00001010, 
8'b11111001, 
8'b00000010, 
8'b11110000, 
8'b00001000, 
8'b00001001, 
8'b00000001, 
8'b11111011, 
8'b00000101, 
8'b11111100, 
8'b00000100, 
8'b00000010, 
8'b00000000, 
8'b00000001, 
8'b11110110, 
8'b00000011, 
8'b11111101, 
8'b00000010, 
8'b00001101, 
8'b00001000, 
8'b11111110, 
8'b11110011, 
8'b00000111, 
8'b11110001, 
8'b11111011, 
8'b11111001, 
8'b11111111, 
8'b00001010, 
8'b11111100, 
8'b00000000, 
8'b00001111, 
8'b11111101, 
8'b11111101, 
8'b11111011, 
8'b11111110, 
8'b00001000, 
8'b11110100, 
8'b11111010, 
8'b11111010, 
8'b11110011, 
8'b11110111, 
8'b11101111, 
8'b11111001, 
8'b11111001, 
8'b11101111, 
8'b00001100, 
8'b11110011, 
8'b00000100, 
8'b11110101, 
8'b11110101, 
8'b00000111, 
8'b00000000, 
8'b11110100, 
8'b00000010, 
8'b11110010, 
8'b00001010, 
8'b00000100, 
8'b11111011, 
8'b11110111, 
8'b11111000, 
8'b00000110, 
8'b11110100, 
8'b00000000, 
8'b00001010, 
8'b00000101, 
8'b00000110, 
8'b11110100, 
8'b00001100, 
8'b00001001, 
8'b00000001, 
8'b00001110, 
8'b00000001, 
8'b11101110, 
8'b00001101, 
8'b00000101, 
8'b00001011, 
8'b11110001, 
8'b11111101, 
8'b00000011, 
8'b11110100, 
8'b11110110, 
8'b11110110, 
8'b11111001, 
8'b00001110, 
8'b00000000, 
8'b00000110, 
8'b00000000, 
8'b00001100, 
8'b00001011, 
8'b11110000, 
8'b11110101, 
8'b00001000, 
8'b11110111, 
8'b11111101, 
8'b11111101, 
8'b00001000, 
8'b00000011, 
8'b11111111, 
8'b11110101, 
8'b00001001, 
8'b11111100, 
8'b00001010, 
8'b00000011, 
8'b00000101, 
8'b11111011, 
8'b00000001, 
8'b00001010, 
8'b11111101, 
8'b11111111, 
8'b11111110, 
8'b11110110, 
8'b00010000, 
8'b00000010, 
8'b11111000, 
8'b11111110, 
8'b00000011, 
8'b11111101, 
8'b11111101, 
8'b00000010, 
8'b00001100, 
8'b00000111, 
8'b00001011, 
8'b00000011, 
8'b11110110, 
8'b00000010, 
8'b11110110, 
8'b11111010, 
8'b11111000, 
8'b00000000, 
8'b00000001, 
8'b00000101, 
8'b00000011, 
8'b00000100, 
8'b11101100, 
8'b11110110, 
8'b11111110, 
8'b00000001, 
8'b00001111, 
8'b00001111, 
8'b11101111, 
8'b11111101, 
8'b00001000, 
8'b00001101, 
8'b11101111, 
8'b11110110, 
8'b00000001, 
8'b00001001, 
8'b11111010, 
8'b11111011, 
8'b11111100, 
8'b11111111, 
8'b00001101, 
8'b00001010, 
8'b11111110, 
8'b11111011, 
8'b00001001, 
8'b00000100, 
8'b00001000, 
8'b11111110, 
8'b11111000, 
8'b11111100, 
8'b11111110, 
8'b11110010, 
8'b00000010, 
8'b11110011, 
8'b00000110, 
8'b11111110, 
8'b11111110, 
8'b00001000, 
8'b00000001, 
8'b11111110, 
8'b00000101, 
8'b00000100, 
8'b00000011, 
8'b00000001, 
8'b00000110, 
8'b11110111, 
8'b00010000, 
8'b00000111, 
8'b11101110, 
8'b00000001, 
8'b11110010, 
8'b11110001, 
8'b11101101, 
8'b11111100, 
8'b11111010, 
8'b11111000, 
8'b00000101, 
8'b00000001, 
8'b11110011, 
8'b00000010, 
8'b11111000, 
8'b11111001, 
8'b11111010, 
8'b11111011, 
8'b11111001, 
8'b00000001, 
8'b11111100, 
8'b00001001, 
8'b11111000, 
8'b00000011, 
8'b00000001, 
8'b00000101, 
8'b00001101, 
8'b00000000, 
8'b11110111, 
8'b11111010, 
8'b00000111, 
8'b00001000, 
8'b11101011, 
8'b00000100, 
8'b00000001, 
8'b11101110, 
8'b00001011, 
8'b11111011, 
8'b00000000, 
8'b11110110, 
8'b00001011, 
8'b00000111, 
8'b11101001, 
8'b00001000, 
8'b00000101, 
8'b00000101, 
8'b00010010, 
8'b00000101, 
8'b00001010, 
8'b11110110, 
8'b00000010, 
8'b11111100, 
8'b00000100, 
8'b00001110, 
8'b00000111, 
8'b11101011, 
8'b00001010, 
8'b11111011, 
8'b00000010, 
8'b11110111, 
8'b11110100, 
8'b00000010, 
8'b00000111, 
8'b00000011, 
8'b11111100, 
8'b11101101, 
8'b00000100, 
8'b00000001, 
8'b00001001, 
8'b00000000, 
8'b00000010, 
8'b00001001, 
8'b00001000, 
8'b11111011, 
8'b00000110, 
8'b11110111, 
8'b11110111, 
8'b11111010, 
8'b00001011, 
8'b11111000, 
8'b11110100, 
8'b00000001, 
8'b00000110, 
8'b00001000, 
8'b11111001, 
8'b11101110, 
8'b11101110, 
8'b00000111, 
8'b00000000, 
8'b00001010, 
8'b00001000, 
8'b00000111, 
8'b00001011, 
8'b11111010, 
8'b11111111, 
8'b00000010, 
8'b00000100, 
8'b00001001, 
8'b00001010, 
8'b00001101, 
8'b11110111, 
8'b00000000, 
8'b00001101, 
8'b00001001, 
8'b00001001, 
8'b11111111, 
8'b11110101, 
8'b11111101, 
8'b11111101, 
8'b11110111, 
8'b11110000, 
8'b00001000, 
8'b00000111, 
8'b00001010, 
8'b00000000, 
8'b11111001, 
8'b11111101, 
8'b11111000, 
8'b00000001, 
8'b00000000, 
8'b00001011, 
8'b00000101, 
8'b11101110, 
8'b11110110, 
8'b11110100, 
8'b11111111, 
8'b11110001, 
8'b11111100, 
8'b11111011, 
8'b00000011, 
8'b00000000, 
8'b00000010, 
8'b11101100, 
8'b11111111, 
8'b00001000, 
8'b00001101, 
8'b11111110, 
8'b11110000, 
8'b00000111, 
8'b11111100, 
8'b00001011, 
8'b11111111, 
8'b11101101, 
8'b11111010, 
8'b00000001, 
8'b11110001, 
8'b11111110, 
8'b00001011, 
8'b11111011, 
8'b11111111, 
8'b00001010, 
8'b00000011, 
8'b11111011, 
8'b00001011, 
8'b11111011, 
8'b00000100, 
8'b00000000, 
8'b11110011, 
8'b00001010, 
8'b11111001, 
8'b00000000, 
8'b00000001, 
8'b11111010, 
8'b11111100, 
8'b00000111, 
8'b00000000, 
8'b00000010, 
8'b00000100, 
8'b11111000, 
8'b00000011, 
8'b11110101, 
8'b11111111, 
8'b11111001, 
8'b11111001, 
8'b11110110, 
8'b00000001, 
8'b00000101, 
8'b00000010, 
8'b11111011, 
8'b11110110, 
8'b00001010, 
8'b11111001, 
8'b00000000, 
8'b00001100, 
8'b00000000, 
8'b11110011, 
8'b00001000, 
8'b11110111, 
8'b00000101, 
8'b00000011, 
8'b00000100, 
8'b00001000, 
8'b11110110, 
8'b00000011, 
8'b11111001, 
8'b11110100, 
8'b00000110, 
8'b11110011, 
8'b00001011, 
8'b00000010, 
8'b11111011, 
8'b11110011, 
8'b11111010, 
8'b00001010, 
8'b11111000, 
8'b00000000, 
8'b11111010, 
8'b00001100, 
8'b11111101, 
8'b00000001, 
8'b00000110, 
8'b11111001, 
8'b11111000, 
8'b00000011, 
8'b00000001, 
8'b11110001, 
8'b00001101, 
8'b11111101, 
8'b00001100, 
8'b00000111, 
8'b00000110, 
8'b11110111, 
8'b11111101, 
8'b11111101, 
8'b11111011, 
8'b11111110, 
8'b00000111, 
8'b11111000, 
8'b00000110, 
8'b00000001, 
8'b00000010, 
8'b00000110, 
8'b00001010, 
8'b00000101, 
8'b11111000, 
8'b00000011, 
8'b11110000, 
8'b00000100, 
8'b11111011, 
8'b00000110, 
8'b11111010, 
8'b11111001, 
8'b00000101, 
8'b11110110, 
8'b11111001, 
8'b11110101, 
8'b00000001, 
8'b11111000, 
8'b00001110, 
8'b11111110, 
8'b11111000, 
8'b11111111, 
8'b00000101, 
8'b00000101, 
8'b00001010, 
8'b11111010, 
8'b11110100, 
8'b00000000, 
8'b11110111, 
8'b11111010, 
8'b11110010, 
8'b00000110, 
8'b00010000, 
8'b00000110, 
8'b00001010, 
8'b11111111, 
8'b11111000, 
8'b00001001, 
8'b11111100, 
8'b00001010, 
8'b11111011, 
8'b00000010, 
8'b11110100, 
8'b00010001, 
8'b00001111, 
8'b11111001, 
8'b11101011, 
8'b00000001, 
8'b11110110, 
8'b00010000, 
8'b11111110, 
8'b11111001, 
8'b00000001, 
8'b11111000, 
8'b11111001, 
8'b11111011, 
8'b11101100, 
8'b00000001, 
8'b11101101, 
8'b11111010, 
8'b00000001, 
8'b00000101, 
8'b11111000, 
8'b11111110, 
8'b00000010, 
8'b11111011, 
8'b11101010, 
8'b11111011, 
8'b00000011, 
8'b00000010, 
8'b00000100, 
8'b00000101, 
8'b11101110, 
8'b11111010, 
8'b00001011, 
8'b11110011, 
8'b11111011, 
8'b00001110, 
8'b11111001, 
8'b00000000, 
8'b11111001, 
8'b00000010, 
8'b11111101, 
8'b11111011, 
8'b00001011, 
8'b11110011, 
8'b11111011, 
8'b00001001, 
8'b00001011, 
8'b11111100, 
8'b00000100, 
8'b11111101, 
8'b11101110, 
8'b11111011, 
8'b00000010, 
8'b11111001, 
8'b11111111, 
8'b11111100, 
8'b11111001, 
8'b00001001, 
8'b11111001, 
8'b11111000, 
8'b00000000, 
8'b11111100, 
8'b00000101, 
8'b11110101, 
8'b00001010, 
8'b00000111, 
8'b00000000, 
8'b11111111, 
8'b11110111, 
8'b11110101, 
8'b11111000, 
8'b11111011, 
8'b11111101, 
8'b00000010, 
8'b00001111, 
8'b11111011, 
8'b11110001, 
8'b00001110, 
8'b11111000, 
8'b11111110, 
8'b00000010, 
8'b00000110, 
8'b11110111, 
8'b11111000, 
8'b11111100, 
8'b00000111, 
8'b11111001, 
8'b00000110, 
8'b00000111, 
8'b11110100, 
8'b00000000, 
8'b00000000, 
8'b11111100, 
8'b11111011, 
8'b00000001, 
8'b11111100, 
8'b00000011, 
8'b00000011, 
8'b11110101, 
8'b11111000, 
8'b00000001, 
8'b00000111, 
8'b11110010, 
8'b11101110, 
8'b11111001, 
8'b11111101, 
8'b11111101, 
8'b11111110, 
8'b11110110, 
8'b00000101, 
8'b00000101, 
8'b11111001, 
8'b00000110, 
8'b11111111, 
8'b11111011, 
8'b00001011, 
8'b11111000, 
8'b11111101, 
8'b11111000, 
8'b00000011, 
8'b00001001, 
8'b11111111, 
8'b00000101, 
8'b11101101, 
8'b00000001, 
8'b11111001, 
8'b11111010, 
8'b00001001, 
8'b11110100, 
8'b00000101, 
8'b11111010, 
8'b00000000, 
8'b00000000, 
8'b11110011, 
8'b11111111, 
8'b00000001, 
8'b11110110, 
8'b00000010, 
8'b00001010, 
8'b11111001, 
8'b00000111, 
8'b11111100, 
8'b00001101, 
8'b11101011, 
8'b11101011, 
8'b00000110, 
8'b11111010, 
8'b00000010, 
8'b11110111, 
8'b11111101, 
8'b00000111, 
8'b00000010, 
8'b11111111, 
8'b00000010, 
8'b11111001, 
8'b00001000, 
8'b11111111, 
8'b11111001, 
8'b00000101, 
8'b11111110, 
8'b00000000, 
8'b00000111, 
8'b11110010, 
8'b11111000, 
8'b11101011, 
8'b00000100, 
8'b11110010, 
8'b00000110, 
8'b00000100, 
8'b11111111, 
8'b11110111, 
8'b11111001, 
8'b00000111, 
8'b11111110, 
8'b11101111, 
8'b00001100, 
8'b11101110, 
8'b11110110, 
8'b11111110, 
8'b00000000, 
8'b11110100, 
8'b11111010, 
8'b11111111, 
8'b11111110, 
8'b11111101, 
8'b11111111, 
8'b11111000, 
8'b00001110, 
8'b11111100, 
8'b00000001, 
8'b00000001, 
8'b11111101, 
8'b00000010, 
8'b00000001, 
8'b11111100, 
8'b11111101, 
8'b00000011, 
8'b00000001, 
8'b00000010, 
8'b00000101, 
8'b11110110, 
8'b00001111, 
8'b11111010, 
8'b00000010, 
8'b11111010, 
8'b00000101, 
8'b11110100, 
8'b11110111, 
8'b11110001, 
8'b11111101, 
8'b11101011, 
8'b11111111, 
8'b11111000, 
8'b11110100, 
8'b11110111, 
8'b11111011, 
8'b11111000, 
8'b00001010, 
8'b11101011, 
8'b00010000, 
8'b11111101, 
8'b11110111, 
8'b11111101, 
8'b11110011, 
8'b00000010, 
8'b00000101, 
8'b11110101, 
8'b00000010, 
8'b11110001, 
8'b00001000, 
8'b11110011, 
8'b00000010, 
8'b11111010, 
8'b11111100, 
8'b00001011, 
8'b00001001, 
8'b11111001, 
8'b00001000, 
8'b00000011, 
8'b00000010, 
8'b00001101, 
8'b00000111, 
8'b11111001, 
8'b11111000, 
8'b00001011, 
8'b00001010, 
8'b00000000, 
8'b00000110, 
8'b00000010, 
8'b00000010, 
8'b11111101, 
8'b00001001, 
8'b11111110, 
8'b00000000, 
8'b00000011, 
8'b00010011, 
8'b11110101, 
8'b11111011, 
8'b00000000, 
8'b00001000, 
8'b00001001, 
8'b11110110, 
8'b11110101, 
8'b00000001, 
8'b00000011, 
8'b00000001, 
8'b00000010, 
8'b00000100, 
8'b00000011, 
8'b00001000, 
8'b11111111, 
8'b00000001, 
8'b00001001, 
8'b11111111, 
8'b11111101, 
8'b00000010, 
8'b11110011, 
8'b00000001, 
8'b00000101, 
8'b11110101, 
8'b00001111, 
8'b11111111, 
8'b00000011, 
8'b11111111, 
8'b11111101, 
8'b11111101, 
8'b00000111, 
8'b00001111, 
8'b00000000, 
8'b00000110, 
8'b00010000, 
8'b11110011, 
8'b00000111, 
8'b00001000, 
8'b11110111, 
8'b00000001, 
8'b00001001, 
8'b00000000, 
8'b00000111, 
8'b11111110, 
8'b00001101, 
8'b00000101, 
8'b11111010, 
8'b11110000, 
8'b11110110, 
8'b00000011, 
8'b00000000, 
8'b11111110, 
8'b00000100, 
8'b00000101, 
8'b00000101, 
8'b11110001, 
8'b00000010, 
8'b00000110, 
8'b11110011, 
8'b11111001, 
8'b11111101, 
8'b00001100, 
8'b00001101, 
8'b11111111, 
8'b00000111, 
8'b11110011, 
8'b11111011, 
8'b11111011, 
8'b11111110, 
8'b00000001, 
8'b11101111, 
8'b00000111, 
8'b11111100, 
8'b11111100, 
8'b11110101, 
8'b00000001, 
8'b11111111, 
8'b00010010, 
8'b11110001, 
8'b00000100, 
8'b00000000, 
8'b11111000, 
8'b11111011, 
8'b00000010, 
8'b11110101, 
8'b11111001, 
8'b11110001, 
8'b11111100, 
8'b00000110, 
8'b00001100, 
8'b11110111, 
8'b11111100, 
8'b00000010, 
8'b00001010, 
8'b11111011, 
8'b11111111, 
8'b11111110, 
8'b00001011, 
8'b11101110, 
8'b00001010, 
8'b11111001, 
8'b11101111, 
8'b11110111, 
8'b00010000, 
8'b11110010, 
8'b11111100, 
8'b11110000, 
8'b00000110, 
8'b00001110, 
8'b00001110, 
8'b11110111, 
8'b00000000, 
8'b11101111, 
8'b00000110, 
8'b11111000, 
8'b00001001, 
8'b00000000, 
8'b00000101, 
8'b11111000, 
8'b11111001, 
8'b11110111, 
8'b00000011, 
8'b00000100, 
8'b00001101, 
8'b00000010, 
8'b11111000, 
8'b11111100, 
8'b11110010, 
8'b00001010, 
8'b00000111, 
8'b11110100, 
8'b11111100, 
8'b11101111, 
8'b00001010, 
8'b11110011, 
8'b00001101, 
8'b11110111, 
8'b00000011, 
8'b00000001, 
8'b00001010, 
8'b11110110, 
8'b11110101, 
8'b00001011, 
8'b11111001, 
8'b00000001, 
8'b11110101, 
8'b00000000, 
8'b11111010, 
8'b00000111, 
8'b11111011, 
8'b11111001, 
8'b11111010, 
8'b00000110, 
8'b11111011, 
8'b11111101, 
8'b00000101, 
8'b00001001, 
8'b11110000, 
8'b00000001, 
8'b00000001, 
8'b11101111, 
8'b11111101, 
8'b00001100, 
8'b00000111, 
8'b11110001, 
8'b00000111, 
8'b11100100, 
8'b11110010, 
8'b11110100, 
8'b00000001, 
8'b11101110, 
8'b11111011, 
8'b00000001, 
8'b11111010, 
8'b00001111, 
8'b00000010, 
8'b00000000, 
8'b00000000, 
8'b00010010, 
8'b11110100, 
8'b11110101, 
8'b00000010, 
8'b00001010, 
8'b00001000, 
8'b00001000, 
8'b11111000, 
8'b11110101, 
8'b00000001, 
8'b11110111, 
8'b00000010, 
8'b00000011, 
8'b00000001, 
8'b11110001, 
8'b11110001, 
8'b11111110, 
8'b11111100, 
8'b11111101, 
8'b11110000, 
8'b00000010, 
8'b11111010, 
8'b11101101, 
8'b11110111, 
8'b00001010, 
8'b11110011, 
8'b00001001, 
8'b00010000, 
8'b00001111, 
8'b11111111, 
8'b11110101, 
8'b00000110, 
8'b11110101, 
8'b11111011, 
8'b00000110, 
8'b11111110, 
8'b11111101, 
8'b11111101, 
8'b00001000
};

localparam logic signed [7:0] dlBiases [9:0] = {
8'b00001010, 
8'b11111111, 
8'b11111111, 
8'b11111100, 
8'b11111100, 
8'b11111110, 
8'b11111110, 
8'b00000100, 
8'b11110100, 
8'b11111110
};

localparam logic signed [7:0] convWeights [0:17] = {
8'b00000111, 
8'b00011110, 
8'b11110000, 
8'b00000101, 
8'b00000000, 
8'b00100000, 
8'b00011001, 
8'b00001100, 
8'b11110001, 
8'b00010110, 
8'b11111010, 
8'b00001101, 
8'b00011111, 
8'b00001010, 
8'b00011000, 
8'b11111111, 
8'b00001011, 
8'b00000111
};

localparam logic signed [7:0] convBiases [1:0] = {
8'b00000000, 
8'b00000000
};
endpackage