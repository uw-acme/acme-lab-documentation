package data12_6;
localparam logic signed [11:0] dlWeights [0:1279] = {
12'b000000010000, 
12'b000000000000, 
12'b111111110011, 
12'b000000000000, 
12'b111111111011, 
12'b000000001000, 
12'b000000000100, 
12'b111111110011, 
12'b000000000010, 
12'b000000001010, 
12'b000000001010, 
12'b111111101111, 
12'b111111100111, 
12'b111111110101, 
12'b000000000110, 
12'b111111111000, 
12'b111111111011, 
12'b111111111110, 
12'b111111111100, 
12'b111111111111, 
12'b000000000111, 
12'b111111110000, 
12'b000000000011, 
12'b000000000101, 
12'b111111111101, 
12'b000000000000, 
12'b111111111011, 
12'b000000000010, 
12'b000000000100, 
12'b000000010000, 
12'b000000100100, 
12'b111111100100, 
12'b111111110000, 
12'b111111101101, 
12'b111111110001, 
12'b000000000111, 
12'b111111111110, 
12'b000000001010, 
12'b111111111011, 
12'b000000001101, 
12'b000000001001, 
12'b111111110111, 
12'b111111111110, 
12'b111111110101, 
12'b000000000000, 
12'b111111111001, 
12'b000000001011, 
12'b111111110110, 
12'b111111111000, 
12'b000000000000, 
12'b000000010111, 
12'b111111110110, 
12'b111111101111, 
12'b111111101010, 
12'b111111110101, 
12'b000000000110, 
12'b111111111110, 
12'b000000001000, 
12'b000000000100, 
12'b000000000110, 
12'b000000001111, 
12'b111111110011, 
12'b000000000100, 
12'b000000000100, 
12'b111111110101, 
12'b000000001110, 
12'b000000001101, 
12'b000000000000, 
12'b000000001011, 
12'b111111111010, 
12'b000000000000, 
12'b000000001101, 
12'b111111110001, 
12'b111111110110, 
12'b111111110101, 
12'b000000000110, 
12'b111111111101, 
12'b000000001011, 
12'b111111110001, 
12'b111111110100, 
12'b111111111011, 
12'b111111111001, 
12'b111111110001, 
12'b000000000110, 
12'b111111110111, 
12'b000000001000, 
12'b000000000000, 
12'b111111110101, 
12'b111111111100, 
12'b111111111000, 
12'b000000000010, 
12'b000000000001, 
12'b111111111001, 
12'b000000000001, 
12'b111111101110, 
12'b111111111100, 
12'b111111110000, 
12'b000000010100, 
12'b111111101111, 
12'b111111101100, 
12'b000000000001, 
12'b000000010011, 
12'b000000000000, 
12'b000000000010, 
12'b111111110110, 
12'b111111111110, 
12'b111111110100, 
12'b111111110101, 
12'b000000000110, 
12'b111111110011, 
12'b000000000001, 
12'b000000001010, 
12'b000000000010, 
12'b000000001000, 
12'b111111110000, 
12'b111111111001, 
12'b111111101111, 
12'b000000000111, 
12'b111111110101, 
12'b000000000100, 
12'b111111110100, 
12'b111111111100, 
12'b000000000001, 
12'b000000000100, 
12'b111111110000, 
12'b111111111011, 
12'b111111110001, 
12'b111111111001, 
12'b000000000000, 
12'b000000000101, 
12'b111111110101, 
12'b111111111011, 
12'b111111111001, 
12'b000000010001, 
12'b111111110100, 
12'b111111101011, 
12'b111111110110, 
12'b000000010100, 
12'b111111111100, 
12'b000000000011, 
12'b111111111111, 
12'b111111111010, 
12'b000000000000, 
12'b000000000011, 
12'b000000001100, 
12'b111111111101, 
12'b111111101111, 
12'b000000001101, 
12'b111111111100, 
12'b000000000100, 
12'b000000000001, 
12'b000000000101, 
12'b000000001001, 
12'b111111111111, 
12'b000000000101, 
12'b111111110110, 
12'b111111001111, 
12'b000000001100, 
12'b111111111101, 
12'b000000000110, 
12'b000000001010, 
12'b111111111100, 
12'b111111101111, 
12'b000000001011, 
12'b000000001101, 
12'b111111111001, 
12'b000000010000, 
12'b111111111100, 
12'b000000000010, 
12'b111111111110, 
12'b000000001001, 
12'b111111111111, 
12'b111111111100, 
12'b111111101010, 
12'b000000000001, 
12'b000000000011, 
12'b111111111010, 
12'b111111111110, 
12'b111111111000, 
12'b000000001001, 
12'b000000001111, 
12'b111111110001, 
12'b111111111110, 
12'b111111111010, 
12'b000000001111, 
12'b111111111111, 
12'b000000001000, 
12'b111111111000, 
12'b000000001100, 
12'b000000000000, 
12'b000000001111, 
12'b111111101001, 
12'b111111110110, 
12'b111111101111, 
12'b111111111111, 
12'b000000000101, 
12'b000000000010, 
12'b000000000110, 
12'b000000001001, 
12'b111111111101, 
12'b000000001101, 
12'b111111101111, 
12'b111111111001, 
12'b111111110111, 
12'b111111111111, 
12'b000000000000, 
12'b000000000000, 
12'b111111111101, 
12'b000000000001, 
12'b111111111001, 
12'b111111111100, 
12'b111111111101, 
12'b111111111101, 
12'b111111110010, 
12'b111111111111, 
12'b000000000001, 
12'b000000001101, 
12'b111111111010, 
12'b000000000000, 
12'b000000000010, 
12'b111111110111, 
12'b111111111100, 
12'b111111110011, 
12'b000000001011, 
12'b111111110011, 
12'b000000001111, 
12'b111111110100, 
12'b000000000001, 
12'b111111111010, 
12'b111111101110, 
12'b000000001010, 
12'b000000001110, 
12'b111111110011, 
12'b000000000100, 
12'b111111111110, 
12'b000000000000, 
12'b111111111001, 
12'b000000001010, 
12'b000000000011, 
12'b000000000011, 
12'b000000000000, 
12'b111111111001, 
12'b000000000101, 
12'b000000000111, 
12'b000000000101, 
12'b111111111010, 
12'b111111110101, 
12'b111111111011, 
12'b000000000111, 
12'b111111110110, 
12'b000000000100, 
12'b000000000100, 
12'b111111111011, 
12'b111111110111, 
12'b111111101111, 
12'b111111111001, 
12'b000000000000, 
12'b000000000000, 
12'b111111101100, 
12'b111111110010, 
12'b111111110000, 
12'b000000000010, 
12'b000000000001, 
12'b000000000101, 
12'b111111101010, 
12'b000000000001, 
12'b000000000111, 
12'b111111110010, 
12'b000000000000, 
12'b111111111110, 
12'b000000000001, 
12'b000000001011, 
12'b000000000011, 
12'b000000000001, 
12'b111111111101, 
12'b111111110011, 
12'b111111110001, 
12'b000000010000, 
12'b111111101110, 
12'b000000000001, 
12'b111111111111, 
12'b000000000000, 
12'b000000000101, 
12'b111111111100, 
12'b000000000010, 
12'b111111111001, 
12'b000000000110, 
12'b111111111111, 
12'b000000001001, 
12'b000000000101, 
12'b111111111001, 
12'b000000000111, 
12'b000000000111, 
12'b000000000000, 
12'b000000000101, 
12'b111111111001, 
12'b111111101100, 
12'b111111111110, 
12'b111111110101, 
12'b111111111011, 
12'b000000000010, 
12'b000000001100, 
12'b000000000011, 
12'b000000000101, 
12'b111111111011, 
12'b000000000010, 
12'b000000000101, 
12'b111111111011, 
12'b000000000110, 
12'b000000001100, 
12'b000000000111, 
12'b000000000100, 
12'b111111111101, 
12'b000000000011, 
12'b000000001001, 
12'b000000000101, 
12'b111111110000, 
12'b000000000001, 
12'b111111111101, 
12'b111111111111, 
12'b000000001000, 
12'b111111101110, 
12'b111111110111, 
12'b000000000110, 
12'b000000001101, 
12'b000000000001, 
12'b000000001101, 
12'b111111101111, 
12'b000000000000, 
12'b000000000111, 
12'b000000010001, 
12'b111111101111, 
12'b111111111010, 
12'b111111101011, 
12'b111111111100, 
12'b000000000110, 
12'b111111110111, 
12'b000000000010, 
12'b111111111010, 
12'b111111110110, 
12'b000000000111, 
12'b111111111010, 
12'b111111111100, 
12'b111111110100, 
12'b000000000010, 
12'b111111111011, 
12'b000000000011, 
12'b111111111001, 
12'b000000001010, 
12'b111111110111, 
12'b000000001010, 
12'b111111111011, 
12'b111111101001, 
12'b000000000011, 
12'b000000001001, 
12'b000000000000, 
12'b000000000001, 
12'b000000000010, 
12'b000000001010, 
12'b111111111001, 
12'b000000000010, 
12'b111111110000, 
12'b000000001000, 
12'b000000001001, 
12'b000000000001, 
12'b111111111011, 
12'b000000000101, 
12'b111111111100, 
12'b000000000100, 
12'b000000000010, 
12'b000000000000, 
12'b000000000001, 
12'b111111110110, 
12'b000000000011, 
12'b111111111101, 
12'b000000000010, 
12'b000000001101, 
12'b000000001000, 
12'b111111111110, 
12'b111111110011, 
12'b000000000111, 
12'b111111110001, 
12'b111111111011, 
12'b111111111001, 
12'b111111111111, 
12'b000000001010, 
12'b111111111100, 
12'b000000000000, 
12'b000000001111, 
12'b111111111101, 
12'b111111111101, 
12'b111111111011, 
12'b111111111110, 
12'b000000001000, 
12'b111111110100, 
12'b111111111010, 
12'b111111111010, 
12'b111111110011, 
12'b111111110111, 
12'b111111101111, 
12'b111111111001, 
12'b111111111001, 
12'b111111101111, 
12'b000000001100, 
12'b111111110011, 
12'b000000000100, 
12'b111111110101, 
12'b111111110101, 
12'b000000000111, 
12'b000000000000, 
12'b111111110100, 
12'b000000000010, 
12'b111111110010, 
12'b000000001010, 
12'b000000000100, 
12'b111111111011, 
12'b111111110111, 
12'b111111111000, 
12'b000000000110, 
12'b111111110100, 
12'b000000000000, 
12'b000000001010, 
12'b000000000101, 
12'b000000000110, 
12'b111111110100, 
12'b000000001100, 
12'b000000001001, 
12'b000000000001, 
12'b000000001110, 
12'b000000000001, 
12'b111111101110, 
12'b000000001101, 
12'b000000000101, 
12'b000000001011, 
12'b111111110001, 
12'b111111111101, 
12'b000000000011, 
12'b111111110100, 
12'b111111110110, 
12'b111111110110, 
12'b111111111001, 
12'b000000001110, 
12'b000000000000, 
12'b000000000110, 
12'b000000000000, 
12'b000000001100, 
12'b000000001011, 
12'b111111110000, 
12'b111111110101, 
12'b000000001000, 
12'b111111110111, 
12'b111111111101, 
12'b111111111101, 
12'b000000001000, 
12'b000000000011, 
12'b111111111111, 
12'b111111110101, 
12'b000000001001, 
12'b111111111100, 
12'b000000001010, 
12'b000000000011, 
12'b000000000101, 
12'b111111111011, 
12'b000000000001, 
12'b000000001010, 
12'b111111111101, 
12'b111111111111, 
12'b111111111110, 
12'b111111110110, 
12'b000000010000, 
12'b000000000010, 
12'b111111111000, 
12'b111111111110, 
12'b000000000011, 
12'b111111111101, 
12'b111111111101, 
12'b000000000010, 
12'b000000001100, 
12'b000000000111, 
12'b000000001011, 
12'b000000000011, 
12'b111111110110, 
12'b000000000010, 
12'b111111110110, 
12'b111111111010, 
12'b111111111000, 
12'b000000000000, 
12'b000000000001, 
12'b000000000101, 
12'b000000000011, 
12'b000000000100, 
12'b111111101100, 
12'b111111110110, 
12'b111111111110, 
12'b000000000001, 
12'b000000001111, 
12'b000000001111, 
12'b111111101111, 
12'b111111111101, 
12'b000000001000, 
12'b000000001101, 
12'b111111101111, 
12'b111111110110, 
12'b000000000001, 
12'b000000001001, 
12'b111111111010, 
12'b111111111011, 
12'b111111111100, 
12'b111111111111, 
12'b000000001101, 
12'b000000001010, 
12'b111111111110, 
12'b111111111011, 
12'b000000001001, 
12'b000000000100, 
12'b000000001000, 
12'b111111111110, 
12'b111111111000, 
12'b111111111100, 
12'b111111111110, 
12'b111111110010, 
12'b000000000010, 
12'b111111110011, 
12'b000000000110, 
12'b111111111110, 
12'b111111111110, 
12'b000000001000, 
12'b000000000001, 
12'b111111111110, 
12'b000000000101, 
12'b000000000100, 
12'b000000000011, 
12'b000000000001, 
12'b000000000110, 
12'b111111110111, 
12'b000000010000, 
12'b000000000111, 
12'b111111101110, 
12'b000000000001, 
12'b111111110010, 
12'b111111110001, 
12'b111111101101, 
12'b111111111100, 
12'b111111111010, 
12'b111111111000, 
12'b000000000101, 
12'b000000000001, 
12'b111111110011, 
12'b000000000010, 
12'b111111111000, 
12'b111111111001, 
12'b111111111010, 
12'b111111111011, 
12'b111111111001, 
12'b000000000001, 
12'b111111111100, 
12'b000000001001, 
12'b111111111000, 
12'b000000000011, 
12'b000000000001, 
12'b000000000101, 
12'b000000001101, 
12'b000000000000, 
12'b111111110111, 
12'b111111111010, 
12'b000000000111, 
12'b000000001000, 
12'b111111101011, 
12'b000000000100, 
12'b000000000001, 
12'b111111101110, 
12'b000000001011, 
12'b111111111011, 
12'b000000000000, 
12'b111111110110, 
12'b000000001011, 
12'b000000000111, 
12'b111111101001, 
12'b000000001000, 
12'b000000000101, 
12'b000000000101, 
12'b000000010010, 
12'b000000000101, 
12'b000000001010, 
12'b111111110110, 
12'b000000000010, 
12'b111111111100, 
12'b000000000100, 
12'b000000001110, 
12'b000000000111, 
12'b111111101011, 
12'b000000001010, 
12'b111111111011, 
12'b000000000010, 
12'b111111110111, 
12'b111111110100, 
12'b000000000010, 
12'b000000000111, 
12'b000000000011, 
12'b111111111100, 
12'b111111101101, 
12'b000000000100, 
12'b000000000001, 
12'b000000001001, 
12'b000000000000, 
12'b000000000010, 
12'b000000001001, 
12'b000000001000, 
12'b111111111011, 
12'b000000000110, 
12'b111111110111, 
12'b111111110111, 
12'b111111111010, 
12'b000000001011, 
12'b111111111000, 
12'b111111110100, 
12'b000000000001, 
12'b000000000110, 
12'b000000001000, 
12'b111111111001, 
12'b111111101110, 
12'b111111101110, 
12'b000000000111, 
12'b000000000000, 
12'b000000001010, 
12'b000000001000, 
12'b000000000111, 
12'b000000001011, 
12'b111111111010, 
12'b111111111111, 
12'b000000000010, 
12'b000000000100, 
12'b000000001001, 
12'b000000001010, 
12'b000000001101, 
12'b111111110111, 
12'b000000000000, 
12'b000000001101, 
12'b000000001001, 
12'b000000001001, 
12'b111111111111, 
12'b111111110101, 
12'b111111111101, 
12'b111111111101, 
12'b111111110111, 
12'b111111110000, 
12'b000000001000, 
12'b000000000111, 
12'b000000001010, 
12'b000000000000, 
12'b111111111001, 
12'b111111111101, 
12'b111111111000, 
12'b000000000001, 
12'b000000000000, 
12'b000000001011, 
12'b000000000101, 
12'b111111101110, 
12'b111111110110, 
12'b111111110100, 
12'b111111111111, 
12'b111111110001, 
12'b111111111100, 
12'b111111111011, 
12'b000000000011, 
12'b000000000000, 
12'b000000000010, 
12'b111111101100, 
12'b111111111111, 
12'b000000001000, 
12'b000000001101, 
12'b111111111110, 
12'b111111110000, 
12'b000000000111, 
12'b111111111100, 
12'b000000001011, 
12'b111111111111, 
12'b111111101101, 
12'b111111111010, 
12'b000000000001, 
12'b111111110001, 
12'b111111111110, 
12'b000000001011, 
12'b111111111011, 
12'b111111111111, 
12'b000000001010, 
12'b000000000011, 
12'b111111111011, 
12'b000000001011, 
12'b111111111011, 
12'b000000000100, 
12'b000000000000, 
12'b111111110011, 
12'b000000001010, 
12'b111111111001, 
12'b000000000000, 
12'b000000000001, 
12'b111111111010, 
12'b111111111100, 
12'b000000000111, 
12'b000000000000, 
12'b000000000010, 
12'b000000000100, 
12'b111111111000, 
12'b000000000011, 
12'b111111110101, 
12'b111111111111, 
12'b111111111001, 
12'b111111111001, 
12'b111111110110, 
12'b000000000001, 
12'b000000000101, 
12'b000000000010, 
12'b111111111011, 
12'b111111110110, 
12'b000000001010, 
12'b111111111001, 
12'b000000000000, 
12'b000000001100, 
12'b000000000000, 
12'b111111110011, 
12'b000000001000, 
12'b111111110111, 
12'b000000000101, 
12'b000000000011, 
12'b000000000100, 
12'b000000001000, 
12'b111111110110, 
12'b000000000011, 
12'b111111111001, 
12'b111111110100, 
12'b000000000110, 
12'b111111110011, 
12'b000000001011, 
12'b000000000010, 
12'b111111111011, 
12'b111111110011, 
12'b111111111010, 
12'b000000001010, 
12'b111111111000, 
12'b000000000000, 
12'b111111111010, 
12'b000000001100, 
12'b111111111101, 
12'b000000000001, 
12'b000000000110, 
12'b111111111001, 
12'b111111111000, 
12'b000000000011, 
12'b000000000001, 
12'b111111110001, 
12'b000000001101, 
12'b111111111101, 
12'b000000001100, 
12'b000000000111, 
12'b000000000110, 
12'b111111110111, 
12'b111111111101, 
12'b111111111101, 
12'b111111111011, 
12'b111111111110, 
12'b000000000111, 
12'b111111111000, 
12'b000000000110, 
12'b000000000001, 
12'b000000000010, 
12'b000000000110, 
12'b000000001010, 
12'b000000000101, 
12'b111111111000, 
12'b000000000011, 
12'b111111110000, 
12'b000000000100, 
12'b111111111011, 
12'b000000000110, 
12'b111111111010, 
12'b111111111001, 
12'b000000000101, 
12'b111111110110, 
12'b111111111001, 
12'b111111110101, 
12'b000000000001, 
12'b111111111000, 
12'b000000001110, 
12'b111111111110, 
12'b111111111000, 
12'b111111111111, 
12'b000000000101, 
12'b000000000101, 
12'b000000001010, 
12'b111111111010, 
12'b111111110100, 
12'b000000000000, 
12'b111111110111, 
12'b111111111010, 
12'b111111110010, 
12'b000000000110, 
12'b000000010000, 
12'b000000000110, 
12'b000000001010, 
12'b111111111111, 
12'b111111111000, 
12'b000000001001, 
12'b111111111100, 
12'b000000001010, 
12'b111111111011, 
12'b000000000010, 
12'b111111110100, 
12'b000000010001, 
12'b000000001111, 
12'b111111111001, 
12'b111111101011, 
12'b000000000001, 
12'b111111110110, 
12'b000000010000, 
12'b111111111110, 
12'b111111111001, 
12'b000000000001, 
12'b111111111000, 
12'b111111111001, 
12'b111111111011, 
12'b111111101100, 
12'b000000000001, 
12'b111111101101, 
12'b111111111010, 
12'b000000000001, 
12'b000000000101, 
12'b111111111000, 
12'b111111111110, 
12'b000000000010, 
12'b111111111011, 
12'b111111101010, 
12'b111111111011, 
12'b000000000011, 
12'b000000000010, 
12'b000000000100, 
12'b000000000101, 
12'b111111101110, 
12'b111111111010, 
12'b000000001011, 
12'b111111110011, 
12'b111111111011, 
12'b000000001110, 
12'b111111111001, 
12'b000000000000, 
12'b111111111001, 
12'b000000000010, 
12'b111111111101, 
12'b111111111011, 
12'b000000001011, 
12'b111111110011, 
12'b111111111011, 
12'b000000001001, 
12'b000000001011, 
12'b111111111100, 
12'b000000000100, 
12'b111111111101, 
12'b111111101110, 
12'b111111111011, 
12'b000000000010, 
12'b111111111001, 
12'b111111111111, 
12'b111111111100, 
12'b111111111001, 
12'b000000001001, 
12'b111111111001, 
12'b111111111000, 
12'b000000000000, 
12'b111111111100, 
12'b000000000101, 
12'b111111110101, 
12'b000000001010, 
12'b000000000111, 
12'b000000000000, 
12'b111111111111, 
12'b111111110111, 
12'b111111110101, 
12'b111111111000, 
12'b111111111011, 
12'b111111111101, 
12'b000000000010, 
12'b000000001111, 
12'b111111111011, 
12'b111111110001, 
12'b000000001110, 
12'b111111111000, 
12'b111111111110, 
12'b000000000010, 
12'b000000000110, 
12'b111111110111, 
12'b111111111000, 
12'b111111111100, 
12'b000000000111, 
12'b111111111001, 
12'b000000000110, 
12'b000000000111, 
12'b111111110100, 
12'b000000000000, 
12'b000000000000, 
12'b111111111100, 
12'b111111111011, 
12'b000000000001, 
12'b111111111100, 
12'b000000000011, 
12'b000000000011, 
12'b111111110101, 
12'b111111111000, 
12'b000000000001, 
12'b000000000111, 
12'b111111110010, 
12'b111111101110, 
12'b111111111001, 
12'b111111111101, 
12'b111111111101, 
12'b111111111110, 
12'b111111110110, 
12'b000000000101, 
12'b000000000101, 
12'b111111111001, 
12'b000000000110, 
12'b111111111111, 
12'b111111111011, 
12'b000000001011, 
12'b111111111000, 
12'b111111111101, 
12'b111111111000, 
12'b000000000011, 
12'b000000001001, 
12'b111111111111, 
12'b000000000101, 
12'b111111101101, 
12'b000000000001, 
12'b111111111001, 
12'b111111111010, 
12'b000000001001, 
12'b111111110100, 
12'b000000000101, 
12'b111111111010, 
12'b000000000000, 
12'b000000000000, 
12'b111111110011, 
12'b111111111111, 
12'b000000000001, 
12'b111111110110, 
12'b000000000010, 
12'b000000001010, 
12'b111111111001, 
12'b000000000111, 
12'b111111111100, 
12'b000000001101, 
12'b111111101011, 
12'b111111101011, 
12'b000000000110, 
12'b111111111010, 
12'b000000000010, 
12'b111111110111, 
12'b111111111101, 
12'b000000000111, 
12'b000000000010, 
12'b111111111111, 
12'b000000000010, 
12'b111111111001, 
12'b000000001000, 
12'b111111111111, 
12'b111111111001, 
12'b000000000101, 
12'b111111111110, 
12'b000000000000, 
12'b000000000111, 
12'b111111110010, 
12'b111111111000, 
12'b111111101011, 
12'b000000000100, 
12'b111111110010, 
12'b000000000110, 
12'b000000000100, 
12'b111111111111, 
12'b111111110111, 
12'b111111111001, 
12'b000000000111, 
12'b111111111110, 
12'b111111101111, 
12'b000000001100, 
12'b111111101110, 
12'b111111110110, 
12'b111111111110, 
12'b000000000000, 
12'b111111110100, 
12'b111111111010, 
12'b111111111111, 
12'b111111111110, 
12'b111111111101, 
12'b111111111111, 
12'b111111111000, 
12'b000000001110, 
12'b111111111100, 
12'b000000000001, 
12'b000000000001, 
12'b111111111101, 
12'b000000000010, 
12'b000000000001, 
12'b111111111100, 
12'b111111111101, 
12'b000000000011, 
12'b000000000001, 
12'b000000000010, 
12'b000000000101, 
12'b111111110110, 
12'b000000001111, 
12'b111111111010, 
12'b000000000010, 
12'b111111111010, 
12'b000000000101, 
12'b111111110100, 
12'b111111110111, 
12'b111111110001, 
12'b111111111101, 
12'b111111101011, 
12'b111111111111, 
12'b111111111000, 
12'b111111110100, 
12'b111111110111, 
12'b111111111011, 
12'b111111111000, 
12'b000000001010, 
12'b111111101011, 
12'b000000010000, 
12'b111111111101, 
12'b111111110111, 
12'b111111111101, 
12'b111111110011, 
12'b000000000010, 
12'b000000000101, 
12'b111111110101, 
12'b000000000010, 
12'b111111110001, 
12'b000000001000, 
12'b111111110011, 
12'b000000000010, 
12'b111111111010, 
12'b111111111100, 
12'b000000001011, 
12'b000000001001, 
12'b111111111001, 
12'b000000001000, 
12'b000000000011, 
12'b000000000010, 
12'b000000001101, 
12'b000000000111, 
12'b111111111001, 
12'b111111111000, 
12'b000000001011, 
12'b000000001010, 
12'b000000000000, 
12'b000000000110, 
12'b000000000010, 
12'b000000000010, 
12'b111111111101, 
12'b000000001001, 
12'b111111111110, 
12'b000000000000, 
12'b000000000011, 
12'b000000010011, 
12'b111111110101, 
12'b111111111011, 
12'b000000000000, 
12'b000000001000, 
12'b000000001001, 
12'b111111110110, 
12'b111111110101, 
12'b000000000001, 
12'b000000000011, 
12'b000000000001, 
12'b000000000010, 
12'b000000000100, 
12'b000000000011, 
12'b000000001000, 
12'b111111111111, 
12'b000000000001, 
12'b000000001001, 
12'b111111111111, 
12'b111111111101, 
12'b000000000010, 
12'b111111110011, 
12'b000000000001, 
12'b000000000101, 
12'b111111110101, 
12'b000000001111, 
12'b111111111111, 
12'b000000000011, 
12'b111111111111, 
12'b111111111101, 
12'b111111111101, 
12'b000000000111, 
12'b000000001111, 
12'b000000000000, 
12'b000000000110, 
12'b000000010000, 
12'b111111110011, 
12'b000000000111, 
12'b000000001000, 
12'b111111110111, 
12'b000000000001, 
12'b000000001001, 
12'b000000000000, 
12'b000000000111, 
12'b111111111110, 
12'b000000001101, 
12'b000000000101, 
12'b111111111010, 
12'b111111110000, 
12'b111111110110, 
12'b000000000011, 
12'b000000000000, 
12'b111111111110, 
12'b000000000100, 
12'b000000000101, 
12'b000000000101, 
12'b111111110001, 
12'b000000000010, 
12'b000000000110, 
12'b111111110011, 
12'b111111111001, 
12'b111111111101, 
12'b000000001100, 
12'b000000001101, 
12'b111111111111, 
12'b000000000111, 
12'b111111110011, 
12'b111111111011, 
12'b111111111011, 
12'b111111111110, 
12'b000000000001, 
12'b111111101111, 
12'b000000000111, 
12'b111111111100, 
12'b111111111100, 
12'b111111110101, 
12'b000000000001, 
12'b111111111111, 
12'b000000010010, 
12'b111111110001, 
12'b000000000100, 
12'b000000000000, 
12'b111111111000, 
12'b111111111011, 
12'b000000000010, 
12'b111111110101, 
12'b111111111001, 
12'b111111110001, 
12'b111111111100, 
12'b000000000110, 
12'b000000001100, 
12'b111111110111, 
12'b111111111100, 
12'b000000000010, 
12'b000000001010, 
12'b111111111011, 
12'b111111111111, 
12'b111111111110, 
12'b000000001011, 
12'b111111101110, 
12'b000000001010, 
12'b111111111001, 
12'b111111101111, 
12'b111111110111, 
12'b000000010000, 
12'b111111110010, 
12'b111111111100, 
12'b111111110000, 
12'b000000000110, 
12'b000000001110, 
12'b000000001110, 
12'b111111110111, 
12'b000000000000, 
12'b111111101111, 
12'b000000000110, 
12'b111111111000, 
12'b000000001001, 
12'b000000000000, 
12'b000000000101, 
12'b111111111000, 
12'b111111111001, 
12'b111111110111, 
12'b000000000011, 
12'b000000000100, 
12'b000000001101, 
12'b000000000010, 
12'b111111111000, 
12'b111111111100, 
12'b111111110010, 
12'b000000001010, 
12'b000000000111, 
12'b111111110100, 
12'b111111111100, 
12'b111111101111, 
12'b000000001010, 
12'b111111110011, 
12'b000000001101, 
12'b111111110111, 
12'b000000000011, 
12'b000000000001, 
12'b000000001010, 
12'b111111110110, 
12'b111111110101, 
12'b000000001011, 
12'b111111111001, 
12'b000000000001, 
12'b111111110101, 
12'b000000000000, 
12'b111111111010, 
12'b000000000111, 
12'b111111111011, 
12'b111111111001, 
12'b111111111010, 
12'b000000000110, 
12'b111111111011, 
12'b111111111101, 
12'b000000000101, 
12'b000000001001, 
12'b111111110000, 
12'b000000000001, 
12'b000000000001, 
12'b111111101111, 
12'b111111111101, 
12'b000000001100, 
12'b000000000111, 
12'b111111110001, 
12'b000000000111, 
12'b111111100100, 
12'b111111110010, 
12'b111111110100, 
12'b000000000001, 
12'b111111101110, 
12'b111111111011, 
12'b000000000001, 
12'b111111111010, 
12'b000000001111, 
12'b000000000010, 
12'b000000000000, 
12'b000000000000, 
12'b000000010010, 
12'b111111110100, 
12'b111111110101, 
12'b000000000010, 
12'b000000001010, 
12'b000000001000, 
12'b000000001000, 
12'b111111111000, 
12'b111111110101, 
12'b000000000001, 
12'b111111110111, 
12'b000000000010, 
12'b000000000011, 
12'b000000000001, 
12'b111111110001, 
12'b111111110001, 
12'b111111111110, 
12'b111111111100, 
12'b111111111101, 
12'b111111110000, 
12'b000000000010, 
12'b111111111010, 
12'b111111101101, 
12'b111111110111, 
12'b000000001010, 
12'b111111110011, 
12'b000000001001, 
12'b000000010000, 
12'b000000001111, 
12'b111111111111, 
12'b111111110101, 
12'b000000000110, 
12'b111111110101, 
12'b111111111011, 
12'b000000000110, 
12'b111111111110, 
12'b111111111101, 
12'b111111111101, 
12'b000000001000 

};
localparam logic signed [11:0] dlBiases [9:0] = {
12'b000000001010, 
12'b111111111111, 
12'b111111111111, 
12'b111111111100, 
12'b111111111100, 
12'b111111111110, 
12'b111111111110, 
12'b000000000100, 
12'b111111110100, 
12'b111111111110 

};
localparam logic signed [11:0] convWeights [0:17] = {
12'b000000000111, 
12'b000000011110, 
12'b111111110000, 
12'b000000000101, 
12'b000000000000, 
12'b000000100000, 
12'b000000011001, 
12'b000000001100, 
12'b111111110001, 
12'b000000010110, 
12'b111111111010, 
12'b000000001101, 
12'b000000011111, 
12'b000000001010, 
12'b000000011000, 
12'b111111111111, 
12'b000000001011, 
12'b000000000111

};
localparam logic signed [11:0] convBiases [1:0] = {
12'b000000000000, 
12'b000000000000

};
endpackage