package data16_10;

localparam logic signed [15:0] convWeights [0:71] = {
16'b0000000010010010,
16'b0000000011111101,
16'b1111111101110100,
16'b1111111101001001,
16'b1111111111101001,
16'b0000000000101100,
16'b1111111101000110,
16'b1111111111000011,
16'b1111111111110101,
16'b1111110110100001,
16'b1111111001111000,
16'b0000000000110000,
16'b1111110110001001,
16'b1111111100111001,
16'b0000000010111111,
16'b0000000000101100,
16'b0000000001001110,
16'b0000000001000000,
16'b0000010001111110,
16'b0000001110010110,
16'b0000000000101110,
16'b0000010000010101,
16'b0000001100011000,
16'b1111111111101101,
16'b1111111111101101,
16'b1111111111101100,
16'b0000000000001101,
16'b1111111111111101,
16'b0000000110110111,
16'b0000000001000111,
16'b0000000101011100,
16'b0000001111101101,
16'b0000001001101010,
16'b0000000101010011,
16'b0000000110101011,
16'b0000000010000010,
16'b0000000000010101,
16'b1111111000110101,
16'b1111111101110011,
16'b1111111100010111,
16'b1111110010000001,
16'b1111110111010000,
16'b1111111011101000,
16'b1111111011110000,
16'b1111111101110100,
16'b0000001001001011,
16'b1111111111001100,
16'b0000000100001111,
16'b0000000000100011,
16'b0000000000101010,
16'b0000001001000000,
16'b0000000000100010,
16'b1111111111100011,
16'b1111111111110111,
16'b0000000001010001,
16'b0000001001001011,
16'b0000000100000010,
16'b0000000000101010,
16'b0000000000101000,
16'b1111111110010010,
16'b1111111111001100,
16'b1111111111100111,
16'b0000000000000000,
16'b0000000001110011,
16'b1111111111010001,
16'b1111111111011010,
16'b0000000100101000,
16'b1111111100110011,
16'b0000000001001000,
16'b0000000000010111,
16'b1111111101111110,
16'b0000000000011011
};

localparam logic signed [15:0] convBiases [7:0] = {
16'b0000000010001111,
16'b0000000010010010,
16'b0000000000000011,
16'b0000000000000001,
16'b0000000010001110,
16'b1111111110101010,
16'b1111111110100101,
16'b0000000000101101 
};

localparam logic signed [15:0] dlWeights [2047:0] = {
16'b0000000000101111, 
16'b0000000010011011, 
16'b1111110001011110, 
16'b0000001101111101, 
16'b0000001011011010, 
16'b0000000010001000, 
16'b0000010000011010, 
16'b0000000001011001, 
16'b1111110110000011, 
16'b0000000101110010, 
16'b1111111110011001, 
16'b1111111100011111, 
16'b0000000100010100, 
16'b0000000000000010, 
16'b0000000101110111, 
16'b0000000010111001, 
16'b1111111111010110, 
16'b0000001000001010, 
16'b1111111010001101, 
16'b1111111101011011, 
16'b0000000010110111, 
16'b1111111101110100, 
16'b1111111001110111, 
16'b0000001101100100, 
16'b1111111111010000, 
16'b0000000011011011, 
16'b1111110101111110, 
16'b1111111110011010, 
16'b0000000010110110, 
16'b0000000010001001, 
16'b1111111010100010, 
16'b0000000000101111, 
16'b0000000100100000, 
16'b0000000011110100, 
16'b1111110100000101, 
16'b1111111000100111, 
16'b0000000011000111, 
16'b0000000000000111, 
16'b0000000111010010, 
16'b0000000001111111, 
16'b0000000011101101, 
16'b0000000100010001, 
16'b1111111001100100, 
16'b1111111110010111, 
16'b0000000001111101, 
16'b1111111011101001, 
16'b1111111111000111, 
16'b0000000110100010, 
16'b0000000011101110, 
16'b0000000010011101, 
16'b1111110110001101, 
16'b1111111100100110, 
16'b0000000010011000, 
16'b1111111110001101, 
16'b0000000110001111, 
16'b0000000011110100, 
16'b0000000000101010, 
16'b0000000001110010, 
16'b1111111001111101, 
16'b1111111011111101, 
16'b0000000010110101, 
16'b0000000101010001, 
16'b0000001011000011, 
16'b0000000001010111, 
16'b1111111111111011, 
16'b0000000011000100, 
16'b1111110101101001, 
16'b1111111000101110, 
16'b1111111111010010, 
16'b1111111110001011, 
16'b0000001000011111, 
16'b0000000011001010, 
16'b0000000000100011, 
16'b0000000101011101, 
16'b1111111010001111, 
16'b1111111001000101, 
16'b0000000000110110, 
16'b0000000111111000, 
16'b0000000010001100, 
16'b0000000100010011, 
16'b0000000101000111, 
16'b0000000100101000, 
16'b0000010101001111, 
16'b0000001010010001, 
16'b0000000010100011, 
16'b0000000001000100, 
16'b1111111111010111, 
16'b0000000010011111, 
16'b0000000010000110, 
16'b0000000010010011, 
16'b0000010110010101, 
16'b0000000110010101, 
16'b0000000100001100, 
16'b0000000010001100, 
16'b0000000001111001, 
16'b0000000011010001, 
16'b0000000001100110, 
16'b0000001011000101, 
16'b1111111111111100, 
16'b1111111110111110, 
16'b0000000011100010, 
16'b0000000000001100, 
16'b0000001100011111, 
16'b0000000101110101, 
16'b0000000011110010, 
16'b0000000001110100, 
16'b1111110110101011, 
16'b1111110101101111, 
16'b1111111101001011, 
16'b1111111100111001, 
16'b0000001100101100, 
16'b0000000100001110, 
16'b0000000001000000, 
16'b0000000110001100, 
16'b0000010011010101, 
16'b0000001010000010, 
16'b0000000001110010, 
16'b0000000010100100, 
16'b0000000000001101, 
16'b0000000100011111, 
16'b0000000100111011, 
16'b0000000011001010, 
16'b0000010010110000, 
16'b0000000111101101, 
16'b0000000010001100, 
16'b1111111101110001, 
16'b1111111101101110, 
16'b0000000010000101, 
16'b0000000000000111, 
16'b0000001001101111, 
16'b0000000111101100, 
16'b1111110101010111, 
16'b1111111110110100, 
16'b1111111101011100, 
16'b0000001001101110, 
16'b0000000011010110, 
16'b1111110010001000, 
16'b0000000001110010, 
16'b0000000000111111, 
16'b0000010100000000, 
16'b0000001111111100, 
16'b0000000111110000, 
16'b1111111000011110, 
16'b0000000001111110, 
16'b1111111011110011, 
16'b1111111101101010, 
16'b1111111010111000, 
16'b1111110110101110, 
16'b1111110100000111, 
16'b1111111011011111, 
16'b1111111000010001, 
16'b0000001011100001, 
16'b0000000111111001, 
16'b0000000101011101, 
16'b1111111100100011, 
16'b1111111001010110, 
16'b1111111011001011, 
16'b0000010010111010, 
16'b1111111110101111, 
16'b0000000100001001, 
16'b0000000011111110, 
16'b1111101000001011, 
16'b1111110101111000, 
16'b0000000000111111, 
16'b0000000011000111, 
16'b1111110100011000, 
16'b1111110011100001, 
16'b1111101110110100, 
16'b0000000111000110, 
16'b1111111111000011, 
16'b1111111110100110, 
16'b0000000011100011, 
16'b0000000011101011, 
16'b0000010101011010, 
16'b0000001111100010, 
16'b1111111010001010, 
16'b0000000011010010, 
16'b0000001010001011, 
16'b0000001101010100, 
16'b0000010010000100, 
16'b0000001111110001, 
16'b0000000000100100, 
16'b1111111000000101, 
16'b0000000000011110, 
16'b0000000101011110, 
16'b1111111101011111, 
16'b1111111011110010, 
16'b1111110100111000, 
16'b1111110111111101, 
16'b0000001010111001, 
16'b1111110011101101, 
16'b1111111110001111, 
16'b1111110111010011, 
16'b1111110111101101, 
16'b1111111011110011, 
16'b0000000010010011, 
16'b0000000000011111, 
16'b1111111001111101, 
16'b1111111010101000, 
16'b1111111000111101, 
16'b1111110100101111, 
16'b1111111000101100, 
16'b1111111100011011, 
16'b0000001110101000, 
16'b0000000111111101, 
16'b1111101101100000, 
16'b0000010111011011, 
16'b1111111001111001, 
16'b0000000000111110, 
16'b0000000111111110, 
16'b0000000010110011, 
16'b1111111111010111, 
16'b0000000011011001, 
16'b0000000010111101, 
16'b0000000001111110, 
16'b0000000000100101, 
16'b0000000100101111, 
16'b0000000001100101, 
16'b0000000001110010, 
16'b1111111110011011, 
16'b0000000011110011, 
16'b0000000000100000, 
16'b1111111110101010, 
16'b0000000001010111, 
16'b0000000110010110, 
16'b0000000010010001, 
16'b1111111111011000, 
16'b1111110001100010, 
16'b1111110010001100, 
16'b0000000111111010, 
16'b1111111111011110, 
16'b0000000001000001, 
16'b0000000000101011, 
16'b0000000000010101, 
16'b1111111011010000, 
16'b0000000000110010, 
16'b0000000010100000, 
16'b0000001000010110, 
16'b0000000011000001, 
16'b0000000100000010, 
16'b0000000101000101, 
16'b0000000010100010, 
16'b0000000010110111, 
16'b1111111100000110, 
16'b0000000001110101, 
16'b0000000100110000, 
16'b0000000010000011, 
16'b0000000100101010, 
16'b0000000000100111, 
16'b0000000110011101, 
16'b0000000111000100, 
16'b1111111010100000, 
16'b0000000110101010, 
16'b1111111110100110, 
16'b0000000011011000, 
16'b0000000101111011, 
16'b0000001100010101, 
16'b0000000110101000, 
16'b1111111101100000, 
16'b1111110101001011, 
16'b1111111101011000, 
16'b0000001000010001, 
16'b0000001001111010, 
16'b0000000101110110, 
16'b0000000111000100, 
16'b1111110110111011, 
16'b1111110001001001, 
16'b0000001000111001, 
16'b0000000101111011, 
16'b1111111101111110, 
16'b1111111000101000, 
16'b0000000100001110, 
16'b1111111011111011, 
16'b1111111101101000, 
16'b1111111000110011, 
16'b0000001000110010, 
16'b0000000010011000, 
16'b1111111100100010, 
16'b0000001000101101, 
16'b0000000010011001, 
16'b1111111101101001, 
16'b0000010000001110, 
16'b0000000111101001, 
16'b0000000100010100, 
16'b0000001101101110, 
16'b0000001011101011, 
16'b1111111111010011, 
16'b0000000110010001, 
16'b0000000011101000, 
16'b1111111101001110, 
16'b1111110101011111, 
16'b0000000100111001, 
16'b0000000011000011, 
16'b0000000100010001, 
16'b1111110111011011, 
16'b0000000010001111, 
16'b1111111000010001, 
16'b0000000100101100, 
16'b1111111011000100, 
16'b0000001100110100, 
16'b0000000111100010, 
16'b0000000011000001, 
16'b0000011000000111, 
16'b0000000111001100, 
16'b1111111101010011, 
16'b0000000111111100, 
16'b1111111110001100, 
16'b1111110000100000, 
16'b1111110100011010, 
16'b1111111101111000, 
16'b1111110100111010, 
16'b0000001011000101, 
16'b0000000110000000, 
16'b0000001000111010, 
16'b1111111101010100, 
16'b1111101101001011, 
16'b1111110011001101, 
16'b0000001000010001, 
16'b1111110000110101, 
16'b0000000111001011, 
16'b0000001001100000, 
16'b1111111001111000, 
16'b1111110110101101, 
16'b1111110110010010, 
16'b1111111101000101, 
16'b1111111011000010, 
16'b0000001001011010, 
16'b1111110111101100, 
16'b0000000100011101, 
16'b1111110110011101, 
16'b1111110110101100, 
16'b1111111011111010, 
16'b1111111101100101, 
16'b0000001101001111, 
16'b0000011010011110, 
16'b0000000011001001, 
16'b0000000000011101, 
16'b0000000011011000, 
16'b0000010011100001, 
16'b0000000100101010, 
16'b0000000011010110, 
16'b0000000000000000, 
16'b1111111111011100, 
16'b0000000011100110, 
16'b0000000000000001, 
16'b0000000110111010, 
16'b0000010001110000, 
16'b0000000000100000, 
16'b0000000010001001, 
16'b1111111100011001, 
16'b0000000000010011, 
16'b0000000100100001, 
16'b0000000010000010, 
16'b1111111110110110, 
16'b1111111000000000, 
16'b0000001101010010, 
16'b0000001011001111, 
16'b1111111011111011, 
16'b1111111011001110, 
16'b0000000010011010, 
16'b1111111111101100, 
16'b0000000111110110, 
16'b0000000011011010, 
16'b1111111101111110, 
16'b0000000000101101, 
16'b1111111110001011, 
16'b1111101001010001, 
16'b0000000110010011, 
16'b0000000001010000, 
16'b0000000100011110, 
16'b0000001110111011, 
16'b0000000011011010, 
16'b0000000101011100, 
16'b1111111111111001, 
16'b1111111101001100, 
16'b0000000001011111, 
16'b0000000101101000, 
16'b0000000001100111, 
16'b0000010001100000, 
16'b0000000100001110, 
16'b0000000100011000, 
16'b1111111110100000, 
16'b1111111111111001, 
16'b0000000100011011, 
16'b1111110100100101, 
16'b0000001000000000, 
16'b1111110110001111, 
16'b0000010100110110, 
16'b0000001010001001, 
16'b1111110110100110, 
16'b1111111101111111, 
16'b0000001111011110, 
16'b1111011111011010, 
16'b1111111001111100, 
16'b1111110000110011, 
16'b1111111110010110, 
16'b1111111110000001, 
16'b1111111011011010, 
16'b0000001000101111, 
16'b1111111101110010, 
16'b1111110000011001, 
16'b0000010000111001, 
16'b0000001111100010, 
16'b0000001010100010, 
16'b0000001101111101, 
16'b1111111000000011, 
16'b1111010101111100, 
16'b0000000111010101, 
16'b0000000000100111, 
16'b1111111111011110, 
16'b1111111001011111, 
16'b0000001000100111, 
16'b0000000111111001, 
16'b1111111110110110, 
16'b1111111010101001, 
16'b1111111011001111, 
16'b0000000100010101, 
16'b1111111101110001, 
16'b1111101101001111, 
16'b0000010110100101, 
16'b0000001110100111, 
16'b0000000100000001, 
16'b0000100001001101, 
16'b1111110110000000, 
16'b0000001010000011, 
16'b0000001101011110, 
16'b0000000010101010, 
16'b1111111100100110, 
16'b0000000010000100, 
16'b0000010000001111, 
16'b0000001101100000, 
16'b0000000110111101, 
16'b1111111001111011, 
16'b1111110111011001, 
16'b1111110101100011, 
16'b0000000011100011, 
16'b1111111101110011, 
16'b1111101001011111, 
16'b0000000100111110, 
16'b0000000000000011, 
16'b1111111110111101, 
16'b0000000111111011, 
16'b0000000110001000, 
16'b1111111101100110, 
16'b0000000011111100, 
16'b0000010010110110, 
16'b0000011101000101, 
16'b1111111111111011, 
16'b0000000110110111, 
16'b1111111011001001, 
16'b1111111011010101, 
16'b0000001010000011, 
16'b0000001110100111, 
16'b0000000100011000, 
16'b0000100010000011, 
16'b1111110011000111, 
16'b0000000101100110, 
16'b0000001000000011, 
16'b0000001101010110, 
16'b0000000111010001, 
16'b0000001100000111, 
16'b0000000110110111, 
16'b0000010101100111, 
16'b1111111111100111, 
16'b0000000001011101, 
16'b1111111100110011, 
16'b0000001111011000, 
16'b1111101100101110, 
16'b1111111101001001, 
16'b1111111100111000, 
16'b1111111110111001, 
16'b1111111111010111, 
16'b0000000010100111, 
16'b1111111110011011, 
16'b0000001010010010, 
16'b1111101001100110, 
16'b0000000000000010, 
16'b1111111111011000, 
16'b0000000010110000, 
16'b1111111110000100, 
16'b1111111010001100, 
16'b1111110111110001, 
16'b1111110101101110, 
16'b1111111110100100, 
16'b1111111111001010, 
16'b1111111100110001, 
16'b0000001000101011, 
16'b0000000111101010, 
16'b1111111010111011, 
16'b0000000100110100, 
16'b0000000000101110, 
16'b0000001101001100, 
16'b0000001001000001, 
16'b1111111000100010, 
16'b1111110011110011, 
16'b0000000010010011, 
16'b1111111101110111, 
16'b1111111110001101, 
16'b0000001101000111, 
16'b1111101110010000, 
16'b1111111101010110, 
16'b1111111101110111, 
16'b1111111101110001, 
16'b0000000000001111, 
16'b0000000010011011, 
16'b1111111110100100, 
16'b0000001001100001, 
16'b1111101010000011, 
16'b0000000010011000, 
16'b1111111111101001, 
16'b1111111110001001, 
16'b1111111110011101, 
16'b0000000101011011, 
16'b0000000010001101, 
16'b0000000010000011, 
16'b0000000100110111, 
16'b0000001000000101, 
16'b1111110011111110, 
16'b1111110110111110, 
16'b0000000011100101, 
16'b0000001101111101, 
16'b0000000010000001, 
16'b0000000000000001, 
16'b0000001110100101, 
16'b0000010001001111, 
16'b1111111011111001, 
16'b0000010101111000, 
16'b1111111001110101, 
16'b0000000000111001, 
16'b0000000001000110, 
16'b0000010001010001, 
16'b0000000111101100, 
16'b0000001010000010, 
16'b1111111001010100, 
16'b0000001100100111, 
16'b0000000111001111, 
16'b0000000001101010, 
16'b0000000011010110, 
16'b0000000101101110, 
16'b1111110110010110, 
16'b1111111010111110, 
16'b1111111011011000, 
16'b0000000111101001, 
16'b1111111111101001, 
16'b1111111101110110, 
16'b0000000001101110, 
16'b1111111100111100, 
16'b0000000001011101, 
16'b1111111110010101, 
16'b1111111010101000, 
16'b0000000010011110, 
16'b0000001001001011, 
16'b0000000000001101, 
16'b0000000011101000, 
16'b1111111100101110, 
16'b1111111100111111, 
16'b1111111101100011, 
16'b1111110011100100, 
16'b0000001001100000, 
16'b1111111100000011, 
16'b0000000010000100, 
16'b1111111100010000, 
16'b0000000110100101, 
16'b0000000001000101, 
16'b1111111110111001, 
16'b0000000100100000, 
16'b0000000101001110, 
16'b1111111010101101, 
16'b1111111111011000, 
16'b0000000010011111, 
16'b0000000100001000, 
16'b0000000101100000, 
16'b0000000011011011, 
16'b1111110011010110, 
16'b1111101011000001, 
16'b1111111011010001, 
16'b1111111000011010, 
16'b0000001010111110, 
16'b0000000110111000, 
16'b1111110011011001, 
16'b1111111101001111, 
16'b0000000000010011, 
16'b0000001000010001, 
16'b0000000101011011, 
16'b1111111111000000, 
16'b0000000100000101, 
16'b1111111110000010, 
16'b0000000011011110, 
16'b0000000100011000, 
16'b0000010001101111, 
16'b1111110100100000, 
16'b1111111101100101, 
16'b0000000000100101, 
16'b1111111010110101, 
16'b1111111001110111, 
16'b1111111101110010, 
16'b1111111111110000, 
16'b0000000011110101, 
16'b0000000011110111, 
16'b0000000000111110, 
16'b1111111100110110, 
16'b0000000000101100, 
16'b1111110101010010, 
16'b1111111110000110, 
16'b1111111011000111, 
16'b1111111111001010, 
16'b0000000001011010, 
16'b1111111101000010, 
16'b0000000000101110, 
16'b0000001001101010, 
16'b0000000100011011, 
16'b0000000000110101, 
16'b0000000110110101, 
16'b1111111011010101, 
16'b1111110101000100, 
16'b0000000011110000, 
16'b0000000010101101, 
16'b0000000000100000, 
16'b1111111000100111, 
16'b1111111111001111, 
16'b0000000000110011, 
16'b1111110110010111, 
16'b0000010101001010, 
16'b1111111111100010, 
16'b1111111111101111, 
16'b1111111101000010, 
16'b1111111000111011, 
16'b1111111010000101, 
16'b1111111100100010, 
16'b0000000010110101, 
16'b1111111111100001, 
16'b1111111111001101, 
16'b1111111100100101, 
16'b1111111110001010, 
16'b1111110110110100, 
16'b1111111100010010, 
16'b1111111110110011, 
16'b0000000011011000, 
16'b0000000010110100, 
16'b1111111101100011, 
16'b0000000110110001, 
16'b1111111111101100, 
16'b1111111000011101, 
16'b0000000010011001, 
16'b0000000111100111, 
16'b1111111011100001, 
16'b1111111011001000, 
16'b0000000000011010, 
16'b1111111101111000, 
16'b1111111110011110, 
16'b1111111110101001, 
16'b0000000000000011, 
16'b0000001011100110, 
16'b1111111010001110, 
16'b0000001110000111, 
16'b1111110110011010, 
16'b1111111101001100, 
16'b0000001110111100, 
16'b1111110111000100, 
16'b0000000010000010, 
16'b0000000101110100, 
16'b1111111101010001, 
16'b0000000001000100, 
16'b0000010110101001, 
16'b0000000001101001, 
16'b0000001000100000, 
16'b1111110001011111, 
16'b1111111010110000, 
16'b0000000110011100, 
16'b0000000010111010, 
16'b0000000100111101, 
16'b1111111111010101, 
16'b0000000001010100, 
16'b0000000010101110, 
16'b1111111010001010, 
16'b0000000001110110, 
16'b0000000010111001, 
16'b1111111101001111, 
16'b1111111111001110, 
16'b0000000110001010, 
16'b0000000001111010, 
16'b0000000101011010, 
16'b1111111101100111, 
16'b0000000101101001, 
16'b0000000011001100, 
16'b1111111001100101, 
16'b0000000100001111, 
16'b0000000001111010, 
16'b0000000001111001, 
16'b0000001000011001, 
16'b1111110011111000, 
16'b0000000001000000, 
16'b0000000110011011, 
16'b1111111100101010, 
16'b0000000110100000, 
16'b0000000000110011, 
16'b0000000000110011, 
16'b0000000110001100, 
16'b1111110100000000, 
16'b1111111111101011, 
16'b0000000110110001, 
16'b0000000100001001, 
16'b0000000001110001, 
16'b0000000010001010, 
16'b0000000010010000, 
16'b1111111111101010, 
16'b0000001010101110, 
16'b1111111111101011, 
16'b1111111101000101, 
16'b1111111111001001, 
16'b0000000011100001, 
16'b1111111111000111, 
16'b0000000110101101, 
16'b0000000000010010, 
16'b0000001100001101, 
16'b0000000111001110, 
16'b0000000000101011, 
16'b0000001100011000, 
16'b1111111011010000, 
16'b1111111110001000, 
16'b0000000011011011, 
16'b0000000101011001, 
16'b0000000010101110, 
16'b1111111011101100, 
16'b0000000101000101, 
16'b0000000011010101, 
16'b0000000001101101, 
16'b0000000001011101, 
16'b0000000000111101, 
16'b0000000100101001, 
16'b0000000101000110, 
16'b1111111011001011, 
16'b0000000000111010, 
16'b0000000011111100, 
16'b0000000001000111, 
16'b1111111110000111, 
16'b0000000010001100, 
16'b0000000010000011, 
16'b0000001110100111, 
16'b0000000001010010, 
16'b1111111111011110, 
16'b0000000000001010, 
16'b1111111111100011, 
16'b0000000000111101, 
16'b0000000001101001, 
16'b1111111110110110, 
16'b0000000111101011, 
16'b1111111110111000, 
16'b1111111110001101, 
16'b1111111111011000, 
16'b0000000101111011, 
16'b1111111101010000, 
16'b0000000010001111, 
16'b0000000000010100, 
16'b0000000011011011, 
16'b1111111100001001, 
16'b0000000101010100, 
16'b0000000100011010, 
16'b1111111110110111, 
16'b0000000000100010, 
16'b0000000001000111, 
16'b0000000101000110, 
16'b0000000101011001, 
16'b1111111101011011, 
16'b0000000010001101, 
16'b0000000100011001, 
16'b0000000010111100, 
16'b0000000001011001, 
16'b0000000001000111, 
16'b1111111000110010, 
16'b1111101111100101, 
16'b1111101100100010, 
16'b1111110110000001, 
16'b1111110100001011, 
16'b1111110111111110, 
16'b0000000010011111, 
16'b1111000010001001, 
16'b0000000010011011, 
16'b0000000011011110, 
16'b1111110001111110, 
16'b1111011001011100, 
16'b1111111111010101, 
16'b0000000011110101, 
16'b1111111001111010, 
16'b0000000001010000, 
16'b1111111011000010, 
16'b0000100101111000, 
16'b1111110110111101, 
16'b0000000101100110, 
16'b0000000001101000, 
16'b1111111101100111, 
16'b1111110101100001, 
16'b1111111111110101, 
16'b1111110010000011, 
16'b1111111101100001, 
16'b0000000010010010, 
16'b1111110010010100, 
16'b1111111101001010, 
16'b1111111111111011, 
16'b1111111110100011, 
16'b0000000001000000, 
16'b1111110110011001, 
16'b1111101101101001, 
16'b1111110100111111, 
16'b1111110101001000, 
16'b0000001100000011, 
16'b0000001110100100, 
16'b1111111111000011, 
16'b1111111100011111, 
16'b1111111000111010, 
16'b1111110001001110, 
16'b1111110000010100, 
16'b1111110010000000, 
16'b0000000111011000, 
16'b1111110110010110, 
16'b0000000001000011, 
16'b0000000010000010, 
16'b1111110011110000, 
16'b0000000110100000, 
16'b1111111110001010, 
16'b1111110011001110, 
16'b0000001000101000, 
16'b0000000001101010, 
16'b1111111110110100, 
16'b0000000001001010, 
16'b1111110110011000, 
16'b1111111101010100, 
16'b0000001011000111, 
16'b1111110110011101, 
16'b1111111111100110, 
16'b1111111111100001, 
16'b0000000010101010, 
16'b1111111110000000, 
16'b1111111011010000, 
16'b1111110001100000, 
16'b1111110111101001, 
16'b1111110011100011, 
16'b0000010100000101, 
16'b1111111111001110, 
16'b1111111110011010, 
16'b1111111110110000, 
16'b1111111001011001, 
16'b1111110100101101, 
16'b1111110111000111, 
16'b1111110011001001, 
16'b0000001000010001, 
16'b0000000100100111, 
16'b0000000010011110, 
16'b0000000010100011, 
16'b1111110101111010, 
16'b0000000010010110, 
16'b0000010001011011, 
16'b1111110010100100, 
16'b0000000010111111, 
16'b0000000000010111, 
16'b1111111110001111, 
16'b0000000001110011, 
16'b1111111000011100, 
16'b0000000100001000, 
16'b0000010010000010, 
16'b1111110011000101, 
16'b1111111111011001, 
16'b0000000001111111, 
16'b0000000000111001, 
16'b1111111111001101, 
16'b1111111000110110, 
16'b1111110011010110, 
16'b1111110011010101, 
16'b1111110010101111, 
16'b0000001010011001, 
16'b0000000110000110, 
16'b0000000001011001, 
16'b0000000001111010, 
16'b1111111001010101, 
16'b1111110010110001, 
16'b1111110001110110, 
16'b1111110100111010, 
16'b0000010010010110, 
16'b1111110111100010, 
16'b0000000100011101, 
16'b1111111101101110, 
16'b1111111000010100, 
16'b0000000010011110, 
16'b0000010100000010, 
16'b1111110101001001, 
16'b0000000000010011, 
16'b1111111110001100, 
16'b1111111101100010, 
16'b0000000000101101, 
16'b1111110100111110, 
16'b1111111111011000, 
16'b0000010000000010, 
16'b1111110000110101, 
16'b0000000000011000, 
16'b0000000011000110, 
16'b0000000000101110, 
16'b0000000000011000, 
16'b0000000101011101, 
16'b0000000101110010, 
16'b1111111001000000, 
16'b0000000001001101, 
16'b0000000001110011, 
16'b0000010111110001, 
16'b0000000001011101, 
16'b0000001101110100, 
16'b0000000010000000, 
16'b0000000001000111, 
16'b1111110111101000, 
16'b1111111111100111, 
16'b0000000000111111, 
16'b0000000011111000, 
16'b1111111110000101, 
16'b0000000101001110, 
16'b1111110111011000, 
16'b1111110110010000, 
16'b1111111110010101, 
16'b0000000000111001, 
16'b0000000001110100, 
16'b0000000000100101, 
16'b0000000100100111, 
16'b1111111110001010, 
16'b0000000101111010, 
16'b0000000010110101, 
16'b1111111000110001, 
16'b1111111011110000, 
16'b0000001001101101, 
16'b0000110011101101, 
16'b0000000100111110, 
16'b1111111101101001, 
16'b1111111000101001, 
16'b1111110011010110, 
16'b0000000100110001, 
16'b0000000101000000, 
16'b0000001000111101, 
16'b1111100100111000, 
16'b1111111110010111, 
16'b1111111010111101, 
16'b1111111111111010, 
16'b1111111010110111, 
16'b1111111100001000, 
16'b0000000000100110, 
16'b1111111011100001, 
16'b1111100011000111, 
16'b0000000010110111, 
16'b1111111011010110, 
16'b0000000000001001, 
16'b1111111001000010, 
16'b0000001100101110, 
16'b0000001000110011, 
16'b1111110010101101, 
16'b1111100101001100, 
16'b0000000001010001, 
16'b1111111110110111, 
16'b0000000001110001, 
16'b1111111001101101, 
16'b0000010011100100, 
16'b0000001111011001, 
16'b1111100110010001, 
16'b1111101111100111, 
16'b0000000001011100, 
16'b1111111111100100, 
16'b0000000000110011, 
16'b1111111010101001, 
16'b1111110100011001, 
16'b1111111110110000, 
16'b0000010011001111, 
16'b1111111100011000, 
16'b1111111011011101, 
16'b1111111100100101, 
16'b0000001010000011, 
16'b0000000110011001, 
16'b0000000100001111, 
16'b0000000001000101, 
16'b0000001011010111, 
16'b0000000111101001, 
16'b0000000101100100, 
16'b0000000101001000, 
16'b0000000101011110, 
16'b0000000101110010, 
16'b0000000001011010, 
16'b0000000011111001, 
16'b0000000010000101, 
16'b0000000001010110, 
16'b1111111111101001, 
16'b0000000100101010, 
16'b0000000100010000, 
16'b0000001010100001, 
16'b0000000001000111, 
16'b0000000001001101, 
16'b0000000011001101, 
16'b0000000010110101, 
16'b0000000100011100, 
16'b1111111110111100, 
16'b0000000101111011, 
16'b1111111011111100, 
16'b1111110100111100, 
16'b1111111011000010, 
16'b1111111011010101, 
16'b1111111111011010, 
16'b0000000010100100, 
16'b0000000001111000, 
16'b0000000001010100, 
16'b1111111101100001, 
16'b0000000100010010, 
16'b0000000100010000, 
16'b0000000101100011, 
16'b0000001101101111, 
16'b0000000011011000, 
16'b0000000010001010, 
16'b0000000000011001, 
16'b0000001010000101, 
16'b0000000000011010, 
16'b0000000010001100, 
16'b0000000000110001, 
16'b1111111101000010, 
16'b0000000010110110, 
16'b0000000010010100, 
16'b0000000011000100, 
16'b0000000110111101, 
16'b1111111111110110, 
16'b0000000101101000, 
16'b0000000010110110, 
16'b0000000001100001, 
16'b0000000011000111, 
16'b1111111100011101, 
16'b0000001001011001, 
16'b0000000100010011, 
16'b1111110000000111, 
16'b1111111110000101, 
16'b1111111110110000, 
16'b1111101100011010, 
16'b0000000001100011, 
16'b1111111010001001, 
16'b0000000011011000, 
16'b1111111010101011, 
16'b1111111010111011, 
16'b1111111110001001, 
16'b0000000011000110, 
16'b0000000000111010, 
16'b1111110110110100, 
16'b0000000011011001, 
16'b0000000111110000, 
16'b1111110110001000, 
16'b1111111010000011, 
16'b0000000001000111, 
16'b1111111101100100, 
16'b1111111111011010, 
16'b0000001010111101, 
16'b1111111111010110, 
16'b0000000011010001, 
16'b1111110011101011, 
16'b1111111010010001, 
16'b0000000101011000, 
16'b0000000101101111, 
16'b0000001001101000, 
16'b0000000001000011, 
16'b1111111111011100, 
16'b0000000100011101, 
16'b0000000001001000, 
16'b0000000000111000, 
16'b0000000001010001, 
16'b0000000001001111, 
16'b0000000011010000, 
16'b0000000011111001, 
16'b0000000001001010, 
16'b1111111111101010, 
16'b1111111001000111, 
16'b1111110110110000, 
16'b1111111110001011, 
16'b0000000110100101, 
16'b0000000000000001, 
16'b0000000001100010, 
16'b0000000100001110, 
16'b0000000110100100, 
16'b1111110111010000, 
16'b1111111011101111, 
16'b0000000100000110, 
16'b0000000111000111, 
16'b1111111111110000, 
16'b0000000111101100, 
16'b0000000000101111, 
16'b0000000101110010, 
16'b1111110100011001, 
16'b1111111010000011, 
16'b0000000001011110, 
16'b1111111100010010, 
16'b1111111011101100, 
16'b0000000010000000, 
16'b0000000000000011, 
16'b0000001011010101, 
16'b1111111101111001, 
16'b0000000001100001, 
16'b0000000101010110, 
16'b0000000010001100, 
16'b1111111011011110, 
16'b0000000110000000, 
16'b0000000001101001, 
16'b0000000100101110, 
16'b1111110111001011, 
16'b1111111100110000, 
16'b0000000010010011, 
16'b1111111010101111, 
16'b1111111010101111, 
16'b0000000010000101, 
16'b0000000100001010, 
16'b0000000001110100, 
16'b0000001110001100, 
16'b0000001000101001, 
16'b0000000101100111, 
16'b0000000011010100, 
16'b1111111111001011, 
16'b0000000010110100, 
16'b0000000110011011, 
16'b0000000111010000, 
16'b0000010000011000, 
16'b0000001010011101, 
16'b0000000001110010, 
16'b1111111111100000, 
16'b0000000000111011, 
16'b0000000100010100, 
16'b0000000010111010, 
16'b0000000000010101, 
16'b1111110001001100, 
16'b1111111110000010, 
16'b0000000100011101, 
16'b0000000010010100, 
16'b1111111001101001, 
16'b1111111100101110, 
16'b0000000101011101, 
16'b0000000101010001, 
16'b1111111010101110, 
16'b0000000101010111, 
16'b0000001001111000, 
16'b0000000111010000, 
16'b1111110111100001, 
16'b0000000010111011, 
16'b0000000101101011, 
16'b0000000011010010, 
16'b0000001110001011, 
16'b0000001010110111, 
16'b0000000110110011, 
16'b1111111111011001, 
16'b0000000000110100, 
16'b0000000001010110, 
16'b0000000100110101, 
16'b0000000100101011, 
16'b0000001101111010, 
16'b0000000110110111, 
16'b0000000010011100, 
16'b0000000000000010, 
16'b0000000001010011, 
16'b0000000011011001, 
16'b0000000000010001, 
16'b0000000001101110, 
16'b1111110100001111, 
16'b1111111011100110, 
16'b0000000100010101, 
16'b1111110110101000, 
16'b1111111101110000, 
16'b0000000010011010, 
16'b1111110110001110, 
16'b0000000000110000, 
16'b1111111001001111, 
16'b1111110011111101, 
16'b0000000001000100, 
16'b1111111100000111, 
16'b1111111110010100, 
16'b0000000001101111, 
16'b1111111111111100, 
16'b1111111011101110, 
16'b1111111010100010, 
16'b0000000011111110, 
16'b1111111101100011, 
16'b1111111110011101, 
16'b1111111011111011, 
16'b0000001000110010, 
16'b0000000111101111, 
16'b0000000010101100, 
16'b0000000000011001, 
16'b0000001010000001, 
16'b0000000101100001, 
16'b1111111101010100, 
16'b1111111100001001, 
16'b0000000000110000, 
16'b1111111110010011, 
16'b0000000101000101, 
16'b1111111001001000, 
16'b0000000010111100, 
16'b0000000100101100, 
16'b1111110011110100, 
16'b1111111011000011, 
16'b0000000101110000, 
16'b0000000010100100, 
16'b0000000011100010, 
16'b1111111001000101, 
16'b0000000101101010, 
16'b0000000101011100, 
16'b1111111111011110, 
16'b1111110110011101, 
16'b0000000001001000, 
16'b0000000001010101, 
16'b0000000011011101, 
16'b0000000010110111, 
16'b0000001001000010, 
16'b0000000010000100, 
16'b1111110110010110, 
16'b0000000010011000, 
16'b0000000010010001, 
16'b0000000101110011, 
16'b0000000100010110, 
16'b0000000011110000, 
16'b0000001000101001, 
16'b0000000110000100, 
16'b0000000100101110, 
16'b0000001100100011, 
16'b0000000001010001, 
16'b0000000011110100, 
16'b1111111110101000, 
16'b1111111001110011, 
16'b0000000101100111, 
16'b0000000001011110, 
16'b1111111110010000, 
16'b0000001011111001, 
16'b1111111111100101, 
16'b0000000100100010, 
16'b0000000001010100, 
16'b1111111111011110, 
16'b1111111110100100, 
16'b0000000010001111, 
16'b0000000001000000, 
16'b0000000011000000, 
16'b1111111111100001, 
16'b0000000101011001, 
16'b0000000100101101, 
16'b0000000111100010, 
16'b1111111111011001, 
16'b0000000010011001, 
16'b0000000011000011, 
16'b0000000000010111, 
16'b0000000000001111, 
16'b0000000110101000, 
16'b0000000110010000, 
16'b0000000100110100, 
16'b1111111111101011, 
16'b0000000010110011, 
16'b0000000001001100, 
16'b1111111101111001, 
16'b0000000101001111, 
16'b0000000101001101, 
16'b0000000011010111, 
16'b0000000010011011, 
16'b1111110010010101, 
16'b1111111001010010, 
16'b0000000111000101, 
16'b0000000001101000, 
16'b0000000010110010, 
16'b0000000011001111, 
16'b0000000011010011, 
16'b1111111011111011, 
16'b1111110010001010, 
16'b1111111100101101, 
16'b0000000111011000, 
16'b1111110101110000, 
16'b0000000010010100, 
16'b0000000100110011, 
16'b0000000111111101, 
16'b0000000111001011, 
16'b0000000000100010, 
16'b0000000101111000, 
16'b0000000001010101, 
16'b1111111110000110, 
16'b0000000011011011, 
16'b0000000100011000, 
16'b0000000010001001, 
16'b0000001000101011, 
16'b1111111011111110, 
16'b0000000100001010, 
16'b0000000011101000, 
16'b0000000000100001, 
16'b0000000011011100, 
16'b0000000111111000, 
16'b1111110111001010, 
16'b0000000100001000, 
16'b0000000111111101, 
16'b1111111110100110, 
16'b1111110110101110, 
16'b1111101110010110, 
16'b0000000000001001, 
16'b0000001010010011, 
16'b1111111011001111, 
16'b0000001000110111, 
16'b0000000010100101, 
16'b0000000101000110, 
16'b1111110110011011, 
16'b0000000100001000, 
16'b1111111010001100, 
16'b1111111111010100, 
16'b0000001101100001, 
16'b1111111100011011, 
16'b0000000111001110, 
16'b0000000110011001, 
16'b0000000000111111, 
16'b0000000001111101, 
16'b0000000011001001, 
16'b0000000001001110, 
16'b0000000000110011, 
16'b1111110101011011, 
16'b1111111111000000, 
16'b0000000001011110, 
16'b1111111010010010, 
16'b1111110110010001, 
16'b1111111111111101, 
16'b0000000010000000, 
16'b0000000001110111, 
16'b0000001100000011, 
16'b0000001000001010, 
16'b0000000000111011, 
16'b1111111110100110, 
16'b0000000001000011, 
16'b0000000010001001, 
16'b0000000110001101, 
16'b1111111110010111, 
16'b0000001011000011, 
16'b0000001011000010, 
16'b0000000001100101, 
16'b1111110101111001, 
16'b0000000000111101, 
16'b1111111101011000, 
16'b0000000011101111, 
16'b0000000001000111, 
16'b1111110110001100, 
16'b0000000100110110, 
16'b0000000100000101, 
16'b1111111100011000, 
16'b0000001011111000, 
16'b1111111110010110, 
16'b0000000001100100, 
16'b0000000100111110, 
16'b1111111101010001, 
16'b0000000100011110, 
16'b0000001000000001, 
16'b0000000111001001, 
16'b0000000100101010, 
16'b1111111111101001, 
16'b1111111011100111, 
16'b0000000010101001, 
16'b1111110100111101, 
16'b1111111101100111, 
16'b0000000011111111, 
16'b0000000000100110, 
16'b0000000001100101, 
16'b1111111111110010, 
16'b1111111001100100, 
16'b1111111111111101, 
16'b1111110110010010, 
16'b0000000001100100, 
16'b0000000100100011, 
16'b0000001101010100, 
16'b1111111011101100, 
16'b0000000000111101, 
16'b1111111111100000, 
16'b0000000100110101, 
16'b0000000100010001, 
16'b1111111000111100, 
16'b0000000101000100, 
16'b1111111111001110, 
16'b0000000011101110, 
16'b1111111110100111, 
16'b1111111111111110, 
16'b0000000010101110, 
16'b0000001000110000, 
16'b1111111000011110, 
16'b0000000100000001, 
16'b0000000001101010, 
16'b0000000000111000, 
16'b0000000010011001, 
16'b0000000000001100, 
16'b0000000010011011, 
16'b1111111000011100, 
16'b1111111011010100, 
16'b0000000010101110, 
16'b1111111111010000, 
16'b0000000001100110, 
16'b0000000011110101, 
16'b1111111110101100, 
16'b0000000011101010, 
16'b1111110110011000, 
16'b1111111011100000, 
16'b0000000010000111, 
16'b0000000010000001, 
16'b0000000100010110, 
16'b0000000010010010, 
16'b0000000010101010, 
16'b0000000011110111, 
16'b0000000111110101, 
16'b1111110100001001, 
16'b0000000001001000, 
16'b0000000010011010, 
16'b1111111110111000, 
16'b0000000010101100, 
16'b0000000001111100, 
16'b0000000100010100, 
16'b0000000100100100, 
16'b1111111000001100, 
16'b0000000001100001, 
16'b0000000010110000, 
16'b0000000000000101, 
16'b0000000011100101, 
16'b1111111000000111, 
16'b0000001101100100, 
16'b0000001101110111, 
16'b0000000111011101, 
16'b0000000000101110, 
16'b0000000001010100, 
16'b1111101000110000, 
16'b0000001010011111, 
16'b0000000111100100, 
16'b1111111110111011, 
16'b1111111001100011, 
16'b1111110101010011, 
16'b1111111101111110, 
16'b0000000001101110, 
16'b0000000100001000, 
16'b1111110101101001, 
16'b1111111110010101, 
16'b1111111001100011, 
16'b1111111000001011, 
16'b0000010001010100, 
16'b0000000111000001, 
16'b0000000001010001, 
16'b1111110111100101, 
16'b0000001001101100, 
16'b0000000111110001, 
16'b1111111110100011, 
16'b1111111000110000, 
16'b0000000010100011, 
16'b1111111111010011, 
16'b1111011111100011, 
16'b0000000111001001, 
16'b1111111100110100, 
16'b0000000110110011, 
16'b1111111010000001, 
16'b1111111100101110, 
16'b1111110100011100, 
16'b1111111110100111, 
16'b0000001110100100, 
16'b1111111100001100, 
16'b1111111100011010, 
16'b0000000100011001, 
16'b1111111011110100, 
16'b1111111100010000, 
16'b0000000110010000, 
16'b0000000010100010, 
16'b1111111110010111, 
16'b0000011000001111, 
16'b1111111101111001, 
16'b1111111111000100, 
16'b0000000110000100, 
16'b0000000011011010, 
16'b0000000011000011, 
16'b0000000101110101, 
16'b1111110000010011, 
16'b0000011110010001, 
16'b0000000000000010, 
16'b0000000010011101, 
16'b1111111001100101, 
16'b1111110101110111, 
16'b0000000101100100, 
16'b0000000010100001, 
16'b1111101001010010, 
16'b1111101101101000, 
16'b1111111011000001, 
16'b1111111100110001, 
16'b0000000111000101, 
16'b0000000001010000, 
16'b0000001110010001, 
16'b0000001010000010, 
16'b1111111011100100, 
16'b0000001111100001, 
16'b0000001001101101, 
16'b0000000011011110, 
16'b0000000000010110, 
16'b1111111101100111, 
16'b1111111010011110, 
16'b1111111011001110, 
16'b0000000110101001, 
16'b1111110110011010, 
16'b0000000000001100, 
16'b0000000010001010, 
16'b1111111111001001, 
16'b0000000010011000, 
16'b1111110010011110, 
16'b1111111111110011, 
16'b1111111111000100, 
16'b0000000000011001, 
16'b1111111111010100, 
16'b1111111111010101, 
16'b0000000000110000, 
16'b1111111111001100, 
16'b1111110100100001, 
16'b0000000011010010, 
16'b1111111110011000, 
16'b0000000001000111, 
16'b0000000010010011, 
16'b0000001010110011, 
16'b1111111100001000, 
16'b1111110100111111, 
16'b0000001010110111, 
16'b0000001000011011, 
16'b1111111101011000, 
16'b0000011100110011, 
16'b1111111001011101, 
16'b0000000101001111, 
16'b0000000100011001, 
16'b0000000001000001, 
16'b1111111110001111, 
16'b1111111111111110, 
16'b1111110101010011, 
16'b0000010110001100, 
16'b0000000001000101, 
16'b0000000011110111, 
16'b0000000000000011, 
16'b0000000010101010, 
16'b1111110110011000, 
16'b0000000011000101, 
16'b0000000001100111, 
16'b0000000011011110, 
16'b0000000011100010, 
16'b0000000010101010, 
16'b0000000011101101, 
16'b0000000011001101, 
16'b1111110011010100, 
16'b1111111110010110, 
16'b0000000010010110, 
16'b0000000001000101, 
16'b0000000001101001, 
16'b1111111101010000, 
16'b1111111111011111, 
16'b0000000001100001, 
16'b1111111111101100, 
16'b1111111111000000, 
16'b1111111111111001, 
16'b0000000000010101, 
16'b0000000010001100, 
16'b0000000001101111, 
16'b1111111111010001, 
16'b0000000000001010, 
16'b1111111100010111, 
16'b0000000000111100, 
16'b1111111111001010, 
16'b0000000000101110, 
16'b0000000000011101, 
16'b0000000010110010, 
16'b0000000000111101, 
16'b1111111111010010, 
16'b1111111100101010, 
16'b1111111101111110, 
16'b0000000000100011, 
16'b0000000001001001, 
16'b1111111110001111, 
16'b1111111101001110, 
16'b0000000000100001, 
16'b1111111110100001, 
16'b1111111110111110, 
16'b1111111100111101, 
16'b0000000001001000, 
16'b0000000010111100, 
16'b0000000010001001, 
16'b1111111111010100, 
16'b0000000001100010, 
16'b1111111101010111, 
16'b0000000000000100, 
16'b0000000001001011, 
16'b0000000000000000, 
16'b1111111101010100, 
16'b0000000000100001, 
16'b1111111100111010, 
16'b0000000001001101, 
16'b1111111111011110, 
16'b0000000010010000, 
16'b0000000000011011, 
16'b0000000000110110, 
16'b1111111101000011, 
16'b1111111111000101, 
16'b1111111101110001, 
16'b0000000010100011, 
16'b1111111110101000, 
16'b0000000000111010, 
16'b1111111101001101, 
16'b1111111100101001, 
16'b1111111111001010, 
16'b1111111110010011, 
16'b1111111101101000, 
16'b1111111110000001, 
16'b1111111100110100, 
16'b1111111101001100, 
16'b1111111111100000, 
16'b0000000001000100, 
16'b1111111101110011, 
16'b1111111101010100, 
16'b1111111101111101, 
16'b1111111110000010, 
16'b1111111110100011, 
16'b0000000000001000, 
16'b0000000001101011, 
16'b1111111101010110, 
16'b0000000010101100, 
16'b1111111111100111, 
16'b1111111100110111, 
16'b1111111101010001, 
16'b1111111101100000, 
16'b0000000001010000, 
16'b0000000001100110, 
16'b1111111100101111, 
16'b0000000001110100, 
16'b1111111101001110, 
16'b1111111111001101, 
16'b0000000001101100, 
16'b0000000001111001, 
16'b1111111101100010, 
16'b1111111100100100, 
16'b0000000000011100, 
16'b0000000001011101, 
16'b1111111110000001, 
16'b1111111110110010, 
16'b0000000001100001, 
16'b1111111110101001, 
16'b1111111101100010, 
16'b1111111110100011, 
16'b1111111101100001, 
16'b0000000010101000, 
16'b1111111101110110, 
16'b0000000000011010, 
16'b0000000010010100, 
16'b0000000001101000, 
16'b0000000000111111, 
16'b0000000010000000, 
16'b1111111101000010, 
16'b1111111110001111, 
16'b0000000010000010, 
16'b1111111101101101, 
16'b0000000001001001, 
16'b1111111100101101, 
16'b1111111101010111, 
16'b1111111111100100, 
16'b0000000001001011, 
16'b0000000010001100, 
16'b1111111101001110, 
16'b1111111111101011, 
16'b1111111101111011, 
16'b0000000001011010, 
16'b1111111111010011, 
16'b1111111111010101, 
16'b0000000010001100, 
16'b1111111111111010, 
16'b1111111100110110, 
16'b1111111100010001, 
16'b1111111111110011, 
16'b0000000001010111, 
16'b0000000001001110, 
16'b1111111110101010, 
16'b1111111111011001, 
16'b0000000000000110, 
16'b1111111111101010, 
16'b0000000110101001, 
16'b1111110101111100, 
16'b1111111111011110, 
16'b1111110101111110, 
16'b0000000000111100, 
16'b0000001100101101, 
16'b1111110000010000, 
16'b1111110010110010, 
16'b1111111100101001, 
16'b1111111111001100, 
16'b0000010000011100, 
16'b1111101101011100, 
16'b1111111010011011, 
16'b1111110001110101, 
16'b0000000110000110, 
16'b1111101100011000, 
16'b0000000001110100, 
16'b0000001000101010, 
16'b0000001010110101, 
16'b1111110110100100, 
16'b0000000010000000, 
16'b1111111101101111, 
16'b1111111100011001, 
16'b0000000010101000, 
16'b0000000001001100, 
16'b1111111110010000, 
16'b1111111011101001, 
16'b0000001010111001, 
16'b0000001001111000, 
16'b0000000100010100, 
16'b0000001000011100, 
16'b1111111101011000, 
16'b1111111011110011, 
16'b0000000110001011, 
16'b0000001010000001, 
16'b1111111011100111, 
16'b0000000001111100, 
16'b0000000110101000, 
16'b1111110100110011, 
16'b0000000110100000, 
16'b1111111101001001, 
16'b0000000101101101, 
16'b0000001011011111, 
16'b0000001010101111, 
16'b0000000011000111, 
16'b0000000100000111, 
16'b1111101010011010, 
16'b0000000001100010, 
16'b0000000111000011, 
16'b0000000010100001, 
16'b1111111111101001, 
16'b0000000000010011, 
16'b0000000000010111, 
16'b1111111000110111, 
16'b1111111101000000, 
16'b1111111101111100, 
16'b0000000001011110, 
16'b1111111111111110, 
16'b1111110111111001, 
16'b0000001000001101, 
16'b0000000010100010, 
16'b1111111111001110, 
16'b0000010101101111, 
16'b0000000000001010, 
16'b1111111011101111, 
16'b1111111111001100, 
16'b1111110000101111, 
16'b0000010000111110, 
16'b0000000111001001, 
16'b0000000101000110, 
16'b1111111010110101, 
16'b1111111101111011, 
16'b1111111010100111, 
16'b0000000010010110, 
16'b1111111100101011, 
16'b1111111000011110, 
16'b1111111100111011, 
16'b0000000111000001, 
16'b0000010111001111, 
16'b1111111110100110, 
16'b0000000011101101, 
16'b1111111101111100, 
16'b1111111011010110, 
16'b0000000010011100, 
16'b0000000000011110, 
16'b0000000001010101, 
16'b1111111100110101, 
16'b0000000000101000, 
16'b1111111101011111, 
16'b1111111110110011, 
16'b1111111010101011, 
16'b1111111111111100, 
16'b1111111100110101, 
16'b1111111101011000, 
16'b1111111111001101, 
16'b0000000000010111, 
16'b0000000111010100, 
16'b0000000101011010, 
16'b1111111000101100, 
16'b0000000000000011, 
16'b0000000010010100, 
16'b0000010000000101, 
16'b0000100001100000, 
16'b1111111001010100, 
16'b0000000100110011, 
16'b0000000111101010, 
16'b0000000101100010, 
16'b1111110001011101, 
16'b0000000001110000, 
16'b0000011101010100, 
16'b0000000101010001, 
16'b0000000011100011, 
16'b0000000001010110, 
16'b1111111101100010, 
16'b1111110111001011, 
16'b0000000010110011, 
16'b0000000001100110, 
16'b1111111111011001, 
16'b0000000000000000, 
16'b1111111101011101, 
16'b0000000000100101, 
16'b0000000000111111, 
16'b1111111010101000, 
16'b0000000000110000, 
16'b1111111111100111, 
16'b1111111101110100, 
16'b1111111101000010, 
16'b1111111101110000, 
16'b0000000011011101, 
16'b0000000101001111, 
16'b1111010011011010, 
16'b1111100011100111, 
16'b0000000100111000, 
16'b1111010000000001, 
16'b1111101011110110, 
16'b0000000011011010, 
16'b1010011100100100, 
16'b0000000001011100, 
16'b1111111001111010, 
16'b1111100010001110, 
16'b1101001100001100, 
16'b0000000000000010, 
16'b0000001001001100, 
16'b1111111111001011, 
16'b0000000011110010, 
16'b1111011110000101, 
16'b0000000011010001, 
16'b1111110011100111, 
16'b0000000001111000, 
16'b1111111110111110, 
16'b0000000000110101, 
16'b0000010101010010, 
16'b1111111110111011, 
16'b0000000001001010, 
16'b1111001010000100, 
16'b1111101110110001, 
16'b0000000000010111, 
16'b0000000000111111, 
16'b0000000010000101, 
16'b1111111111111100, 
16'b0000000001001101, 
16'b0000000101110010, 
16'b1111001101010000, 
16'b1111101111011110, 
16'b0000000000001110, 
16'b1111110011101010, 
16'b1111111000000111, 
16'b0000000010010111, 
16'b0000000100110011, 
16'b0000000011001010, 
16'b1111010011111000, 
16'b1111101011100000, 
16'b1111111111010111, 
16'b0000010100011011, 
16'b0000010001001001, 
16'b0000000001111110, 
16'b0000000000101001, 
16'b0000000000001111, 
16'b1111010101101011, 
16'b1111110011011100, 
16'b0000000101001101, 
16'b0000001101011010, 
16'b0000001001101100, 
16'b0000000011100111, 
16'b0000000100000101, 
16'b0000000000101010, 
16'b1111000110001011, 
16'b1111101101010111, 
16'b0000000000100010, 
16'b1111111011011110, 
16'b1111100110010001, 
16'b0000000001100100, 
16'b0000000000101010, 
16'b0000000100000000, 
16'b1111011111111010, 
16'b1111110001110011, 
16'b0000000001010111, 
16'b1111101111110011, 
16'b0000000000110000, 
16'b1111111110011101, 
16'b0000000000000000, 
16'b0000000100101000, 
16'b1111100110111100, 
16'b1111110000110111, 
16'b1111111111101001, 
16'b1111100110101110, 
16'b1111100110111000, 
16'b0000000011110101, 
16'b0000000010000100, 
16'b0000000011011010, 
16'b0000010001000011, 
16'b0000000110111000, 
16'b0000000001010011, 
16'b1111111110101101, 
16'b0000000001001001, 
16'b0000000000111001, 
16'b1111111111010111, 
16'b0000000100011000, 
16'b0000010011001110, 
16'b0000001011101001, 
16'b1111111110001111, 
16'b0000000010100001, 
16'b0000000001110011, 
16'b0000000010000011, 
16'b1111111110111010, 
16'b0000000010101000, 
16'b1111101001011111, 
16'b0000000000110000, 
16'b0000000000111100, 
16'b1111111010010010, 
16'b1111011101010111, 
16'b1111111111011000, 
16'b0000000011011110, 
16'b1111111111010100, 
16'b1111100001000000, 
16'b1111101111101001, 
16'b1111111111000111, 
16'b1111111100001001, 
16'b1111011111110011, 
16'b0000000011110001, 
16'b0000000000000101, 
16'b1111111111010101, 
16'b0000010100011010, 
16'b0000001100100110, 
16'b0000000001111110, 
16'b1111111101101010, 
16'b0000000010110010, 
16'b0000000001111111, 
16'b1111111110110110, 
16'b1111111111010101, 
16'b0000010000111011, 
16'b0000001000011010, 
16'b1111111110101001, 
16'b1111111101111001, 
16'b0000000010111000, 
16'b0000000011110101, 
16'b1111111001000010, 
16'b0000000100100110, 
16'b1111110011110011, 
16'b0000000001111000, 
16'b0000000011010110, 
16'b0000001110011010, 
16'b1111110001001010, 
16'b1111111100100001, 
16'b0000000101001000, 
16'b0000000011110000, 
16'b1111111001010011, 
16'b0000000001001111, 
16'b0000001010010100, 
16'b1111111100010100, 
16'b1111111001111001, 
16'b1111111010111111, 
16'b0000000001011111, 
16'b0000000010000100, 
16'b1111111101001010, 
16'b0000001001111110, 
16'b0000000011000000, 
16'b0000000000101011, 
16'b0000010001000000, 
16'b0000000011111010, 
16'b0000000100000000, 
16'b0000000100110100, 
16'b0000000000011001, 
16'b1111110011001011, 
16'b1111110100110010, 
16'b1111110110000111, 
16'b1111101110110100, 
16'b0000000110010010, 
16'b0000000011010110, 
16'b0000000111100101, 
16'b1111111100011000, 
16'b1111111001010111, 
16'b0000000010110110, 
16'b0000001110101101, 
16'b0000010000100011, 
16'b0000000000000110, 
16'b0000000101100101, 
16'b0000000100010000, 
16'b1111111100111010, 
16'b1111110111011111, 
16'b0000000000001000, 
16'b1111110100111111, 
16'b0000000111010100, 
16'b0000000110101101, 
16'b1111111101001001, 
16'b1111111110101011, 
16'b1111111101101100, 
16'b0000000101000010, 
16'b0000000011100110, 
16'b0000001011011101, 
16'b0000001111101101, 
16'b0000000100001011, 
16'b0000000010000000, 
16'b0000000111101010, 
16'b0000000110101000, 
16'b0000000101111001, 
16'b0000000100011110, 
16'b0000000111101110, 
16'b1111110110110110, 
16'b0000000101100100, 
16'b1111111110001110, 
16'b0000000101101010, 
16'b0000000001101011, 
16'b1111111000011111, 
16'b0000000000011101, 
16'b1111111010101101, 
16'b1111100101011111, 
16'b0000000101011000, 
16'b0000000001001101, 
16'b1111111110000110, 
16'b1111111111001101, 
16'b0000000110000100, 
16'b1111111111001110, 
16'b0000000001101100, 
16'b1111101100011101, 
16'b0000000001111001, 
16'b0000000001110100, 
16'b0000000011000011, 
16'b0000000110000110, 
16'b1111111101011100, 
16'b0000000000001100, 
16'b1111111101101110, 
16'b0000000000111101, 
16'b0000000010011101, 
16'b1111111111111010, 
16'b1111111110100101, 
16'b0000000110001011, 
16'b1111111011100001, 
16'b0000000010111100, 
16'b0000000001100011, 
16'b1111111110111100, 
16'b1111111111011111, 
16'b1111111111100010, 
16'b1111111111010001, 
16'b1111111011001001, 
16'b0000000001010111, 
16'b0000000000100010, 
16'b1111111011111011, 
16'b0000000010000100, 
16'b1111111101010111, 
16'b0000000100100100, 
16'b0000000010110111, 
16'b0000000100010000, 
16'b0000001110100000, 
16'b0000001000000001, 
16'b0000001011101011, 
16'b0000010001011001, 
16'b1111111110111011, 
16'b0000000011001111, 
16'b0000000000101000, 
16'b0000000010101100, 
16'b0000000000100000, 
16'b1111111110010100, 
16'b0000000000110001, 
16'b0000000011000111, 
16'b1111111100110101, 
16'b1111111111110000, 
16'b0000000000010110, 
16'b0000001000010001, 
16'b1111111100011011, 
16'b0000000100000111, 
16'b0000000010100101, 
16'b0000000001111001, 
16'b0000000000101000
};

localparam logic signed [15:0] dlBiases [15:0] = {
16'b0000000101010101, 
16'b0000000100000001, 
16'b0000000001111011, 
16'b0000000001000100, 
16'b1111111101111111, 
16'b0000000011101101, 
16'b1111111110110100, 
16'b0000000011100000, 
16'b0000000110001111, 
16'b0000000101001101, 
16'b0000000011011101, 
16'b0000000010010010, 
16'b1111111111011110, 
16'b0000000010010000, 
16'b0000000011100110, 
16'b0000000001111111
};

endpackage