package data14_5;

localparam logic signed [13:0] dlWeights [0:1279] = {
14'b00000010000011, 
14'b00000000000101, 
14'b11111110011100, 
14'b00000000000011, 
14'b11111111011110, 
14'b00000001000100, 
14'b00000000100000, 
14'b11111110011010, 
14'b00000000010111, 
14'b00000001010101, 
14'b00000001010110, 
14'b11111101111011, 
14'b11111100111101, 
14'b11111110101001, 
14'b00000000110001, 
14'b11111111000010, 
14'b11111111011001, 
14'b11111111110000, 
14'b11111111100110, 
14'b11111111111110, 
14'b00000000111101, 
14'b11111110000101, 
14'b00000000011011, 
14'b00000000101001, 
14'b11111111101111, 
14'b00000000000010, 
14'b11111111011110, 
14'b00000000010001, 
14'b00000000100001, 
14'b00000010000001, 
14'b00000100100101, 
14'b11111100100101, 
14'b11111110000011, 
14'b11111101101010, 
14'b11111110001000, 
14'b00000000111110, 
14'b11111111110010, 
14'b00000001010011, 
14'b11111111011011, 
14'b00000001101001, 
14'b00000001001111, 
14'b11111110111010, 
14'b11111111110111, 
14'b11111110101001, 
14'b00000000000010, 
14'b11111111001111, 
14'b00000001011001, 
14'b11111110110011, 
14'b11111111000110, 
14'b00000000000101, 
14'b00000010111010, 
14'b11111110110110, 
14'b11111101111100, 
14'b11111101010100, 
14'b11111110101101, 
14'b00000000110001, 
14'b11111111110100, 
14'b00000001000001, 
14'b00000000100000, 
14'b00000000110100, 
14'b00000001111100, 
14'b11111110011010, 
14'b00000000100001, 
14'b00000000100010, 
14'b11111110101001, 
14'b00000001110100, 
14'b00000001101101, 
14'b00000000000001, 
14'b00000001011001, 
14'b11111111010111, 
14'b00000000000001, 
14'b00000001101011, 
14'b11111110001111, 
14'b11111110110001, 
14'b11111110101110, 
14'b00000000110010, 
14'b11111111101011, 
14'b00000001011010, 
14'b11111110001000, 
14'b11111110100011, 
14'b11111111011001, 
14'b11111111001010, 
14'b11111110001100, 
14'b00000000110101, 
14'b11111110111011, 
14'b00000001000100, 
14'b00000000000000, 
14'b11111110101001, 
14'b11111111100011, 
14'b11111111000111, 
14'b00000000010010, 
14'b00000000001000, 
14'b11111111001001, 
14'b00000000001110, 
14'b11111101110000, 
14'b11111111100101, 
14'b11111110000101, 
14'b00000010100000, 
14'b11111101111011, 
14'b11111101100101, 
14'b00000000001010, 
14'b00000010011000, 
14'b00000000000010, 
14'b00000000010001, 
14'b11111110110011, 
14'b11111111110011, 
14'b11111110100100, 
14'b11111110101010, 
14'b00000000110111, 
14'b11111110011100, 
14'b00000000001110, 
14'b00000001010101, 
14'b00000000010001, 
14'b00000001000001, 
14'b11111110000001, 
14'b11111111001100, 
14'b11111101111001, 
14'b00000000111000, 
14'b11111110101011, 
14'b00000000100000, 
14'b11111110100000, 
14'b11111111100011, 
14'b00000000001000, 
14'b00000000100110, 
14'b11111110000111, 
14'b11111111011110, 
14'b11111110001001, 
14'b11111111001100, 
14'b00000000000001, 
14'b00000000101010, 
14'b11111110101101, 
14'b11111111011111, 
14'b11111111001010, 
14'b00000010001111, 
14'b11111110100110, 
14'b11111101011100, 
14'b11111110110100, 
14'b00000010100010, 
14'b11111111100100, 
14'b00000000011000, 
14'b11111111111001, 
14'b11111111010111, 
14'b00000000000111, 
14'b00000000011000, 
14'b00000001100111, 
14'b11111111101011, 
14'b11111101111001, 
14'b00000001101001, 
14'b11111111100100, 
14'b00000000100011, 
14'b00000000001010, 
14'b00000000101010, 
14'b00000001001010, 
14'b11111111111010, 
14'b00000000101001, 
14'b11111110110101, 
14'b11111001111111, 
14'b00000001100110, 
14'b11111111101001, 
14'b00000000110011, 
14'b00000001010001, 
14'b11111111100010, 
14'b11111101111011, 
14'b00000001011110, 
14'b00000001101110, 
14'b11111111001001, 
14'b00000010000001, 
14'b11111111100010, 
14'b00000000010101, 
14'b11111111110110, 
14'b00000001001011, 
14'b11111111111000, 
14'b11111111100010, 
14'b11111101010001, 
14'b00000000001001, 
14'b00000000011100, 
14'b11111111010101, 
14'b11111111110010, 
14'b11111111000110, 
14'b00000001001011, 
14'b00000001111000, 
14'b11111110001000, 
14'b11111111110111, 
14'b11111111010001, 
14'b00000001111001, 
14'b11111111111011, 
14'b00000001000111, 
14'b11111111000111, 
14'b00000001100101, 
14'b00000000000011, 
14'b00000001111000, 
14'b11111101001110, 
14'b11111110110101, 
14'b11111101111000, 
14'b11111111111100, 
14'b00000000101110, 
14'b00000000010101, 
14'b00000000110101, 
14'b00000001001111, 
14'b11111111101001, 
14'b00000001101000, 
14'b11111101111010, 
14'b11111111001001, 
14'b11111110111010, 
14'b11111111111111, 
14'b00000000000101, 
14'b00000000000001, 
14'b11111111101111, 
14'b00000000001010, 
14'b11111111001100, 
14'b11111111100010, 
14'b11111111101010, 
14'b11111111101001, 
14'b11111110010110, 
14'b11111111111000, 
14'b00000000001101, 
14'b00000001101010, 
14'b11111111010001, 
14'b00000000000111, 
14'b00000000010110, 
14'b11111110111011, 
14'b11111111100110, 
14'b11111110011101, 
14'b00000001011111, 
14'b11111110011011, 
14'b00000001111010, 
14'b11111110100100, 
14'b00000000001001, 
14'b11111111010101, 
14'b11111101110111, 
14'b00000001010001, 
14'b00000001110101, 
14'b11111110011111, 
14'b00000000100011, 
14'b11111111110100, 
14'b00000000000111, 
14'b11111111001010, 
14'b00000001010001, 
14'b00000000011111, 
14'b00000000011001, 
14'b00000000000001, 
14'b11111111001010, 
14'b00000000101010, 
14'b00000000111101, 
14'b00000000101000, 
14'b11111111010110, 
14'b11111110101011, 
14'b11111111011111, 
14'b00000000111100, 
14'b11111110110100, 
14'b00000000100110, 
14'b00000000100011, 
14'b11111111011001, 
14'b11111110111111, 
14'b11111101111010, 
14'b11111111001011, 
14'b00000000000101, 
14'b00000000000000, 
14'b11111101100101, 
14'b11111110010111, 
14'b11111110000000, 
14'b00000000010110, 
14'b00000000001111, 
14'b00000000101101, 
14'b11111101010101, 
14'b00000000001011, 
14'b00000000111000, 
14'b11111110010111, 
14'b00000000000100, 
14'b11111111110011, 
14'b00000000001111, 
14'b00000001011110, 
14'b00000000011010, 
14'b00000000001110, 
14'b11111111101110, 
14'b11111110011000, 
14'b11111110001110, 
14'b00000010000111, 
14'b11111101110010, 
14'b00000000001010, 
14'b11111111111010, 
14'b00000000000100, 
14'b00000000101101, 
14'b11111111100101, 
14'b00000000010001, 
14'b11111111001000, 
14'b00000000110100, 
14'b11111111111111, 
14'b00000001001000, 
14'b00000000101110, 
14'b11111111001000, 
14'b00000000111011, 
14'b00000000111011, 
14'b00000000000010, 
14'b00000000101101, 
14'b11111111001111, 
14'b11111101100100, 
14'b11111111110110, 
14'b11111110101000, 
14'b11111111011101, 
14'b00000000010011, 
14'b00000001100110, 
14'b00000000011000, 
14'b00000000101111, 
14'b11111111011100, 
14'b00000000010100, 
14'b00000000101010, 
14'b11111111011110, 
14'b00000000110011, 
14'b00000001100111, 
14'b00000000111111, 
14'b00000000100110, 
14'b11111111101100, 
14'b00000000011000, 
14'b00000001001011, 
14'b00000000101010, 
14'b11111110000110, 
14'b00000000001001, 
14'b11111111101010, 
14'b11111111111101, 
14'b00000001000010, 
14'b11111101110110, 
14'b11111110111001, 
14'b00000000110110, 
14'b00000001101110, 
14'b00000000001001, 
14'b00000001101111, 
14'b11111101111100, 
14'b00000000000100, 
14'b00000000111101, 
14'b00000010001110, 
14'b11111101111000, 
14'b11111111010100, 
14'b11111101011101, 
14'b11111111100000, 
14'b00000000110011, 
14'b11111110111111, 
14'b00000000010110, 
14'b11111111010011, 
14'b11111110110100, 
14'b00000000111100, 
14'b11111111010100, 
14'b11111111100111, 
14'b11111110100000, 
14'b00000000010011, 
14'b11111111011100, 
14'b00000000011110, 
14'b11111111001011, 
14'b00000001010001, 
14'b11111110111001, 
14'b00000001010001, 
14'b11111111011010, 
14'b11111101001101, 
14'b00000000011001, 
14'b00000001001101, 
14'b00000000000101, 
14'b00000000001101, 
14'b00000000010000, 
14'b00000001010010, 
14'b11111111001110, 
14'b00000000010111, 
14'b11111110000011, 
14'b00000001000000, 
14'b00000001001000, 
14'b00000000001001, 
14'b11111111011110, 
14'b00000000101001, 
14'b11111111100001, 
14'b00000000100010, 
14'b00000000010001, 
14'b00000000000000, 
14'b00000000001100, 
14'b11111110110011, 
14'b00000000011000, 
14'b11111111101001, 
14'b00000000010011, 
14'b00000001101010, 
14'b00000001000101, 
14'b11111111110100, 
14'b11111110011010, 
14'b00000000111001, 
14'b11111110001010, 
14'b11111111011111, 
14'b11111111001111, 
14'b11111111111101, 
14'b00000001010111, 
14'b11111111100101, 
14'b00000000000001, 
14'b00000001111100, 
14'b11111111101000, 
14'b11111111101000, 
14'b11111111011110, 
14'b11111111110110, 
14'b00000001000010, 
14'b11111110100100, 
14'b11111111010011, 
14'b11111111010101, 
14'b11111110011101, 
14'b11111110111100, 
14'b11111101111010, 
14'b11111111001011, 
14'b11111111001110, 
14'b11111101111111, 
14'b00000001100011, 
14'b11111110011111, 
14'b00000000100011, 
14'b11111110101011, 
14'b11111110101100, 
14'b00000000111101, 
14'b00000000000001, 
14'b11111110100101, 
14'b00000000010111, 
14'b11111110010111, 
14'b00000001010010, 
14'b00000000100100, 
14'b11111111011010, 
14'b11111110111101, 
14'b11111111000001, 
14'b00000000110011, 
14'b11111110100000, 
14'b00000000000101, 
14'b00000001010010, 
14'b00000000101100, 
14'b00000000110110, 
14'b11111110100110, 
14'b00000001100111, 
14'b00000001001110, 
14'b00000000001100, 
14'b00000001110100, 
14'b00000000001110, 
14'b11111101110011, 
14'b00000001101100, 
14'b00000000101001, 
14'b00000001011001, 
14'b11111110001110, 
14'b11111111101001, 
14'b00000000011100, 
14'b11111110100111, 
14'b11111110110010, 
14'b11111110110111, 
14'b11111111001011, 
14'b00000001110101, 
14'b00000000000110, 
14'b00000000110100, 
14'b00000000000110, 
14'b00000001100001, 
14'b00000001011100, 
14'b11111110000111, 
14'b11111110101100, 
14'b00000001000110, 
14'b11111110111101, 
14'b11111111101100, 
14'b11111111101100, 
14'b00000001000001, 
14'b00000000011000, 
14'b11111111111011, 
14'b11111110101010, 
14'b00000001001111, 
14'b11111111100101, 
14'b00000001010111, 
14'b00000000011110, 
14'b00000000101010, 
14'b11111111011111, 
14'b00000000001000, 
14'b00000001010111, 
14'b11111111101110, 
14'b11111111111010, 
14'b11111111110100, 
14'b11111110110011, 
14'b00000010000000, 
14'b00000000010011, 
14'b11111111000010, 
14'b11111111110101, 
14'b00000000011100, 
14'b11111111101001, 
14'b11111111101000, 
14'b00000000010010, 
14'b00000001100101, 
14'b00000000111000, 
14'b00000001011011, 
14'b00000000011111, 
14'b11111110110100, 
14'b00000000010100, 
14'b11111110110100, 
14'b11111111010101, 
14'b11111111000010, 
14'b00000000000000, 
14'b00000000001011, 
14'b00000000101011, 
14'b00000000011001, 
14'b00000000100000, 
14'b11111101100111, 
14'b11111110110000, 
14'b11111111110000, 
14'b00000000001110, 
14'b00000001111011, 
14'b00000001111000, 
14'b11111101111001, 
14'b11111111101111, 
14'b00000001000010, 
14'b00000001101011, 
14'b11111101111001, 
14'b11111110110100, 
14'b00000000001110, 
14'b00000001001011, 
14'b11111111010001, 
14'b11111111011101, 
14'b11111111100100, 
14'b11111111111010, 
14'b00000001101011, 
14'b00000001010100, 
14'b11111111110110, 
14'b11111111011011, 
14'b00000001001011, 
14'b00000000100100, 
14'b00000001000101, 
14'b11111111110011, 
14'b11111111000011, 
14'b11111111100011, 
14'b11111111110010, 
14'b11111110010100, 
14'b00000000010110, 
14'b11111110011000, 
14'b00000000110011, 
14'b11111111110000, 
14'b11111111110010, 
14'b00000001000001, 
14'b00000000001001, 
14'b11111111110101, 
14'b00000000101011, 
14'b00000000100001, 
14'b00000000011011, 
14'b00000000001101, 
14'b00000000110000, 
14'b11111110111110, 
14'b00000010000001, 
14'b00000000111111, 
14'b11111101110100, 
14'b00000000001001, 
14'b11111110010000, 
14'b11111110001100, 
14'b11111101101011, 
14'b11111111100101, 
14'b11111111010101, 
14'b11111111000001, 
14'b00000000101101, 
14'b00000000001000, 
14'b11111110011111, 
14'b00000000010100, 
14'b11111111000011, 
14'b11111111001000, 
14'b11111111010000, 
14'b11111111011110, 
14'b11111111001100, 
14'b00000000001000, 
14'b11111111100100, 
14'b00000001001011, 
14'b11111111000000, 
14'b00000000011011, 
14'b00000000001100, 
14'b00000000101100, 
14'b00000001101100, 
14'b00000000000000, 
14'b11111110111010, 
14'b11111111010000, 
14'b00000000111001, 
14'b00000001000111, 
14'b11111101011110, 
14'b00000000100110, 
14'b00000000001001, 
14'b11111101110101, 
14'b00000001011010, 
14'b11111111011000, 
14'b00000000000010, 
14'b11111110110111, 
14'b00000001011000, 
14'b00000000111110, 
14'b11111101001101, 
14'b00000001000111, 
14'b00000000101111, 
14'b00000000101100, 
14'b00000010010100, 
14'b00000000101001, 
14'b00000001010001, 
14'b11111110110001, 
14'b00000000010010, 
14'b11111111100010, 
14'b00000000100010, 
14'b00000001110110, 
14'b00000000111011, 
14'b11111101011101, 
14'b00000001010011, 
14'b11111111011011, 
14'b00000000010110, 
14'b11111110111110, 
14'b11111110100100, 
14'b00000000010001, 
14'b00000000111100, 
14'b00000000011110, 
14'b11111111100011, 
14'b11111101101100, 
14'b00000000100101, 
14'b00000000001101, 
14'b00000001001010, 
14'b00000000000011, 
14'b00000000010001, 
14'b00000001001110, 
14'b00000001000100, 
14'b11111111011011, 
14'b00000000110111, 
14'b11111110111110, 
14'b11111110111111, 
14'b11111111010100, 
14'b00000001011001, 
14'b11111111000011, 
14'b11111110100111, 
14'b00000000001110, 
14'b00000000110111, 
14'b00000001000100, 
14'b11111111001110, 
14'b11111101110111, 
14'b11111101110011, 
14'b00000000111101, 
14'b00000000000111, 
14'b00000001010111, 
14'b00000001000110, 
14'b00000000111011, 
14'b00000001011100, 
14'b11111111010011, 
14'b11111111111000, 
14'b00000000010110, 
14'b00000000100101, 
14'b00000001001110, 
14'b00000001010111, 
14'b00000001101000, 
14'b11111110111100, 
14'b00000000000000, 
14'b00000001101010, 
14'b00000001001101, 
14'b00000001001000, 
14'b11111111111001, 
14'b11111110101111, 
14'b11111111101010, 
14'b11111111101101, 
14'b11111110111100, 
14'b11111110000010, 
14'b00000001000011, 
14'b00000000111100, 
14'b00000001010000, 
14'b00000000000001, 
14'b11111111001111, 
14'b11111111101011, 
14'b11111111000011, 
14'b00000000001111, 
14'b00000000000001, 
14'b00000001011110, 
14'b00000000101001, 
14'b11111101110001, 
14'b11111110110111, 
14'b11111110100101, 
14'b11111111111100, 
14'b11111110001100, 
14'b11111111100111, 
14'b11111111011010, 
14'b00000000011011, 
14'b00000000000100, 
14'b00000000010001, 
14'b11111101100110, 
14'b11111111111010, 
14'b00000001000101, 
14'b00000001101100, 
14'b11111111110101, 
14'b11111110000111, 
14'b00000000111100, 
14'b11111111100011, 
14'b00000001011010, 
14'b11111111111101, 
14'b11111101101111, 
14'b11111111010000, 
14'b00000000001011, 
14'b11111110001001, 
14'b11111111110101, 
14'b00000001011010, 
14'b11111111011010, 
14'b11111111111010, 
14'b00000001010111, 
14'b00000000011101, 
14'b11111111011011, 
14'b00000001011100, 
14'b11111111011100, 
14'b00000000100110, 
14'b00000000000110, 
14'b11111110011101, 
14'b00000001010000, 
14'b11111111001101, 
14'b00000000000100, 
14'b00000000001010, 
14'b11111111010011, 
14'b11111111100110, 
14'b00000000111000, 
14'b00000000000001, 
14'b00000000010110, 
14'b00000000100110, 
14'b11111111000111, 
14'b00000000011101, 
14'b11111110101011, 
14'b11111111111101, 
14'b11111111001101, 
14'b11111111001010, 
14'b11111110110010, 
14'b00000000001100, 
14'b00000000101010, 
14'b00000000010111, 
14'b11111111011000, 
14'b11111110110101, 
14'b00000001010100, 
14'b11111111001111, 
14'b00000000000000, 
14'b00000001100111, 
14'b00000000000010, 
14'b11111110011001, 
14'b00000001000110, 
14'b11111110111001, 
14'b00000000101110, 
14'b00000000011111, 
14'b00000000100000, 
14'b00000001000011, 
14'b11111110110000, 
14'b00000000011001, 
14'b11111111001100, 
14'b11111110100010, 
14'b00000000110111, 
14'b11111110011101, 
14'b00000001011010, 
14'b00000000010001, 
14'b11111111011100, 
14'b11111110011001, 
14'b11111111010011, 
14'b00000001010100, 
14'b11111111000001, 
14'b00000000000101, 
14'b11111111010100, 
14'b00000001100000, 
14'b11111111101111, 
14'b00000000001001, 
14'b00000000110000, 
14'b11111111001101, 
14'b11111111000110, 
14'b00000000011000, 
14'b00000000001100, 
14'b11111110001010, 
14'b00000001101101, 
14'b11111111101001, 
14'b00000001100101, 
14'b00000000111000, 
14'b00000000110010, 
14'b11111110111000, 
14'b11111111101000, 
14'b11111111101000, 
14'b11111111011100, 
14'b11111111110101, 
14'b00000000111000, 
14'b11111111000001, 
14'b00000000110011, 
14'b00000000001011, 
14'b00000000010001, 
14'b00000000110100, 
14'b00000001010000, 
14'b00000000101010, 
14'b11111111000100, 
14'b00000000011101, 
14'b11111110000111, 
14'b00000000100010, 
14'b11111111011010, 
14'b00000000110001, 
14'b11111111010010, 
14'b11111111001001, 
14'b00000000101010, 
14'b11111110110001, 
14'b11111111001111, 
14'b11111110101001, 
14'b00000000001110, 
14'b11111111000110, 
14'b00000001110011, 
14'b11111111110100, 
14'b11111111000100, 
14'b11111111111110, 
14'b00000000101001, 
14'b00000000101000, 
14'b00000001010111, 
14'b11111111010111, 
14'b11111110100000, 
14'b00000000000110, 
14'b11111110111101, 
14'b11111111010111, 
14'b11111110010000, 
14'b00000000110110, 
14'b00000010000110, 
14'b00000000110011, 
14'b00000001010011, 
14'b11111111111100, 
14'b11111111000110, 
14'b00000001001000, 
14'b11111111100001, 
14'b00000001010001, 
14'b11111111011001, 
14'b00000000010111, 
14'b11111110100011, 
14'b00000010001100, 
14'b00000001111001, 
14'b11111111001001, 
14'b11111101011100, 
14'b00000000001011, 
14'b11111110110001, 
14'b00000010000001, 
14'b11111111110000, 
14'b11111111001101, 
14'b00000000001101, 
14'b11111111000110, 
14'b11111111001010, 
14'b11111111011101, 
14'b11111101100111, 
14'b00000000001111, 
14'b11111101101010, 
14'b11111111010101, 
14'b00000000001101, 
14'b00000000101110, 
14'b11111111000111, 
14'b11111111110111, 
14'b00000000010100, 
14'b11111111011011, 
14'b11111101010100, 
14'b11111111011010, 
14'b00000000011010, 
14'b00000000010010, 
14'b00000000100101, 
14'b00000000101000, 
14'b11111101110111, 
14'b11111111010000, 
14'b00000001011000, 
14'b11111110011100, 
14'b11111111011100, 
14'b00000001110111, 
14'b11111111001100, 
14'b00000000000011, 
14'b11111111001110, 
14'b00000000010000, 
14'b11111111101011, 
14'b11111111011100, 
14'b00000001011111, 
14'b11111110011111, 
14'b11111111011100, 
14'b00000001001001, 
14'b00000001011101, 
14'b11111111100101, 
14'b00000000100001, 
14'b11111111101100, 
14'b11111101110100, 
14'b11111111011110, 
14'b00000000010010, 
14'b11111111001110, 
14'b11111111111100, 
14'b11111111100000, 
14'b11111111001110, 
14'b00000001001101, 
14'b11111111001110, 
14'b11111111000000, 
14'b00000000000110, 
14'b11111111100000, 
14'b00000000101000, 
14'b11111110101100, 
14'b00000001010000, 
14'b00000000111111, 
14'b00000000000101, 
14'b11111111111101, 
14'b11111110111000, 
14'b11111110101011, 
14'b11111111000110, 
14'b11111111011011, 
14'b11111111101111, 
14'b00000000010100, 
14'b00000001111001, 
14'b11111111011101, 
14'b11111110001110, 
14'b00000001110101, 
14'b11111111000110, 
14'b11111111110010, 
14'b00000000010001, 
14'b00000000110101, 
14'b11111110111110, 
14'b11111111000100, 
14'b11111111100110, 
14'b00000000111011, 
14'b11111111001110, 
14'b00000000110010, 
14'b00000000111010, 
14'b11111110100110, 
14'b00000000000011, 
14'b00000000000001, 
14'b11111111100110, 
14'b11111111011001, 
14'b00000000001011, 
14'b11111111100111, 
14'b00000000011100, 
14'b00000000011011, 
14'b11111110101001, 
14'b11111111000100, 
14'b00000000001110, 
14'b00000000111100, 
14'b11111110010000, 
14'b11111101110011, 
14'b11111111001110, 
14'b11111111101001, 
14'b11111111101111, 
14'b11111111110110, 
14'b11111110110110, 
14'b00000000101011, 
14'b00000000101111, 
14'b11111111001110, 
14'b00000000110110, 
14'b11111111111000, 
14'b11111111011101, 
14'b00000001011000, 
14'b11111111000011, 
14'b11111111101101, 
14'b11111111000011, 
14'b00000000011001, 
14'b00000001001000, 
14'b11111111111100, 
14'b00000000101101, 
14'b11111101101110, 
14'b00000000001101, 
14'b11111111001011, 
14'b11111111010110, 
14'b00000001001101, 
14'b11111110100011, 
14'b00000000101010, 
14'b11111111010111, 
14'b00000000000010, 
14'b00000000000010, 
14'b11111110011001, 
14'b11111111111001, 
14'b00000000001111, 
14'b11111110110110, 
14'b00000000010000, 
14'b00000001010000, 
14'b11111111001000, 
14'b00000000111100, 
14'b11111111100011, 
14'b00000001101111, 
14'b11111101011111, 
14'b11111101011000, 
14'b00000000110001, 
14'b11111111010010, 
14'b00000000010101, 
14'b11111110111011, 
14'b11111111101011, 
14'b00000000111011, 
14'b00000000010001, 
14'b11111111111100, 
14'b00000000010000, 
14'b11111111001001, 
14'b00000001000101, 
14'b11111111111101, 
14'b11111111001110, 
14'b00000000101000, 
14'b11111111110001, 
14'b00000000000111, 
14'b00000000111110, 
14'b11111110010011, 
14'b11111111000000, 
14'b11111101011110, 
14'b00000000100000, 
14'b11111110010010, 
14'b00000000110000, 
14'b00000000100111, 
14'b11111111111111, 
14'b11111110111111, 
14'b11111111001011, 
14'b00000000111001, 
14'b11111111110100, 
14'b11111101111110, 
14'b00000001100101, 
14'b11111101110001, 
14'b11111110110011, 
14'b11111111110000, 
14'b00000000000000, 
14'b11111110100100, 
14'b11111111010110, 
14'b11111111111110, 
14'b11111111110110, 
14'b11111111101000, 
14'b11111111111010, 
14'b11111111000101, 
14'b00000001110001, 
14'b11111111100010, 
14'b00000000001110, 
14'b00000000001110, 
14'b11111111101100, 
14'b00000000010100, 
14'b00000000001011, 
14'b11111111100111, 
14'b11111111101001, 
14'b00000000011011, 
14'b00000000001101, 
14'b00000000010110, 
14'b00000000101011, 
14'b11111110110100, 
14'b00000001111100, 
14'b11111111010000, 
14'b00000000010000, 
14'b11111111010100, 
14'b00000000101001, 
14'b11111110100111, 
14'b11111110111001, 
14'b11111110001110, 
14'b11111111101010, 
14'b11111101011001, 
14'b11111111111011, 
14'b11111111000111, 
14'b11111110100100, 
14'b11111110111100, 
14'b11111111011111, 
14'b11111111000100, 
14'b00000001010100, 
14'b11111101011110, 
14'b00000010000100, 
14'b11111111101011, 
14'b11111110111101, 
14'b11111111101010, 
14'b11111110011101, 
14'b00000000010010, 
14'b00000000101100, 
14'b11111110101011, 
14'b00000000010111, 
14'b11111110001001, 
14'b00000001000010, 
14'b11111110011111, 
14'b00000000010111, 
14'b11111111010001, 
14'b11111111100001, 
14'b00000001011001, 
14'b00000001001001, 
14'b11111111001100, 
14'b00000001000111, 
14'b00000000011100, 
14'b00000000010011, 
14'b00000001101101, 
14'b00000000111110, 
14'b11111111001000, 
14'b11111111000000, 
14'b00000001011100, 
14'b00000001010101, 
14'b00000000000111, 
14'b00000000110000, 
14'b00000000010111, 
14'b00000000010110, 
14'b11111111101100, 
14'b00000001001111, 
14'b11111111110000, 
14'b00000000000001, 
14'b00000000011110, 
14'b00000010011001, 
14'b11111110101011, 
14'b11111111011101, 
14'b00000000000011, 
14'b00000001000000, 
14'b00000001001111, 
14'b11111110110001, 
14'b11111110101100, 
14'b00000000001010, 
14'b00000000011100, 
14'b00000000001010, 
14'b00000000010000, 
14'b00000000100100, 
14'b00000000011101, 
14'b00000001000010, 
14'b11111111111100, 
14'b00000000001011, 
14'b00000001001000, 
14'b11111111111011, 
14'b11111111101000, 
14'b00000000010000, 
14'b11111110011001, 
14'b00000000001100, 
14'b00000000101100, 
14'b11111110101110, 
14'b00000001111101, 
14'b11111111111000, 
14'b00000000011111, 
14'b11111111111010, 
14'b11111111101101, 
14'b11111111101001, 
14'b00000000111011, 
14'b00000001111110, 
14'b00000000000000, 
14'b00000000110000, 
14'b00000010000001, 
14'b11111110011110, 
14'b00000000111100, 
14'b00000001000001, 
14'b11111110111101, 
14'b00000000001111, 
14'b00000001001110, 
14'b00000000000111, 
14'b00000000111010, 
14'b11111111110111, 
14'b00000001101110, 
14'b00000000101111, 
14'b11111111010001, 
14'b11111110000111, 
14'b11111110110111, 
14'b00000000011001, 
14'b00000000000111, 
14'b11111111110000, 
14'b00000000100011, 
14'b00000000101101, 
14'b00000000101010, 
14'b11111110001100, 
14'b00000000010111, 
14'b00000000110100, 
14'b11111110011011, 
14'b11111111001011, 
14'b11111111101110, 
14'b00000001100100, 
14'b00000001101010, 
14'b11111111111110, 
14'b00000000111010, 
14'b11111110011010, 
14'b11111111011010, 
14'b11111111011110, 
14'b11111111110010, 
14'b00000000001001, 
14'b11111101111000, 
14'b00000000111011, 
14'b11111111100101, 
14'b11111111100100, 
14'b11111110101000, 
14'b00000000001110, 
14'b11111111111011, 
14'b00000010010111, 
14'b11111110001011, 
14'b00000000100000, 
14'b00000000000011, 
14'b11111111000010, 
14'b11111111011001, 
14'b00000000010100, 
14'b11111110101011, 
14'b11111111001110, 
14'b11111110001111, 
14'b11111111100011, 
14'b00000000110111, 
14'b00000001100110, 
14'b11111110111101, 
14'b11111111100110, 
14'b00000000010011, 
14'b00000001010010, 
14'b11111111011110, 
14'b11111111111110, 
14'b11111111110101, 
14'b00000001011000, 
14'b11111101110111, 
14'b00000001010101, 
14'b11111111001000, 
14'b11111101111100, 
14'b11111110111100, 
14'b00000010000101, 
14'b11111110010111, 
14'b11111111100010, 
14'b11111110000001, 
14'b00000000110001, 
14'b00000001110000, 
14'b00000001110110, 
14'b11111110111110, 
14'b00000000000110, 
14'b11111101111001, 
14'b00000000110110, 
14'b11111111000010, 
14'b00000001001011, 
14'b00000000000010, 
14'b00000000101000, 
14'b11111111000001, 
14'b11111111001101, 
14'b11111110111011, 
14'b00000000011001, 
14'b00000000100011, 
14'b00000001101111, 
14'b00000000010001, 
14'b11111111000010, 
14'b11111111100001, 
14'b11111110010010, 
14'b00000001010101, 
14'b00000000111011, 
14'b11111110100010, 
14'b11111111100111, 
14'b11111101111001, 
14'b00000001010101, 
14'b11111110011001, 
14'b00000001101000, 
14'b11111110111111, 
14'b00000000011000, 
14'b00000000001101, 
14'b00000001010000, 
14'b11111110110111, 
14'b11111110101111, 
14'b00000001011010, 
14'b11111111001101, 
14'b00000000001010, 
14'b11111110101010, 
14'b00000000000110, 
14'b11111111010000, 
14'b00000000111010, 
14'b11111111011010, 
14'b11111111001101, 
14'b11111111010000, 
14'b00000000110010, 
14'b11111111011001, 
14'b11111111101010, 
14'b00000000101000, 
14'b00000001001101, 
14'b11111110000101, 
14'b00000000001001, 
14'b00000000001101, 
14'b11111101111100, 
14'b11111111101100, 
14'b00000001100010, 
14'b00000000111010, 
14'b11111110001110, 
14'b00000000111101, 
14'b11111100100010, 
14'b11111110010111, 
14'b11111110100101, 
14'b00000000001000, 
14'b11111101110101, 
14'b11111111011100, 
14'b00000000001001, 
14'b11111111010000, 
14'b00000001111111, 
14'b00000000010000, 
14'b00000000000101, 
14'b00000000000000, 
14'b00000010010110, 
14'b11111110100111, 
14'b11111110101111, 
14'b00000000010111, 
14'b00000001010100, 
14'b00000001000000, 
14'b00000001000001, 
14'b11111111000101, 
14'b11111110101111, 
14'b00000000001111, 
14'b11111110111010, 
14'b00000000010101, 
14'b00000000011111, 
14'b00000000001010, 
14'b11111110001011, 
14'b11111110001010, 
14'b11111111110010, 
14'b11111111100011, 
14'b11111111101101, 
14'b11111110000010, 
14'b00000000010101, 
14'b11111111010100, 
14'b11111101101010, 
14'b11111110111101, 
14'b00000001010111, 
14'b11111110011110, 
14'b00000001001001, 
14'b00000010000001, 
14'b00000001111110, 
14'b11111111111100, 
14'b11111110101011, 
14'b00000000110111, 
14'b11111110101100, 
14'b11111111011100, 
14'b00000000110011, 
14'b11111111110010, 
14'b11111111101111, 
14'b11111111101101, 
14'b00000001000001 
};

localparam logic signed [13:0] dlBiases [9:0] = {
14'b00000001010101, 
14'b11111111111111, 
14'b11111111111111, 
14'b11111111100010, 
14'b11111111100000, 
14'b11111111110101, 
14'b11111111110100, 
14'b00000000100111, 
14'b11111110100011, 
14'b11111111110101
};

localparam logic signed [13:0] convWeights [0:17] = {
14'b00000000111001, 
14'b00000011110110, 
14'b11111110000101, 
14'b00000000101111, 
14'b00000000000111, 
14'b00000100000110, 
14'b00000011001111, 
14'b00000001100110, 
14'b11111110001011, 
14'b00000010110010, 
14'b11111111010011, 
14'b00000001101011, 
14'b00000011111110, 
14'b00000001010001, 
14'b00000011000100, 
14'b11111111111010, 
14'b00000001011101, 
14'b00000000111010
};

localparam logic signed [13:0] convBiases [1:0] = {
14'b00000000000000, 
14'b00000000000000 
};





endpackage