package data6_3;

localparam logic signed [5:0] dlWeights [0:1279] = {
6'b000010, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b000001, 
6'b000001, 
6'b111101, 
6'b111100, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000010, 
6'b000100, 
6'b111100, 
6'b111110, 
6'b111101, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b000001, 
6'b000001, 
6'b111110, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b000010, 
6'b111110, 
6'b111101, 
6'b111101, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b000001, 
6'b000001, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b111110, 
6'b111110, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b111110, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b111110, 
6'b000001, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111101, 
6'b111111, 
6'b111110, 
6'b000010, 
6'b111101, 
6'b111101, 
6'b000000, 
6'b000010, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111110, 
6'b111110, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b000001, 
6'b111110, 
6'b111111, 
6'b111101, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b000010, 
6'b111110, 
6'b111101, 
6'b111110, 
6'b000010, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b111101, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b111001, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b111101, 
6'b000001, 
6'b000001, 
6'b111111, 
6'b000010, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b111101, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b000001, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b000001, 
6'b111101, 
6'b111110, 
6'b111101, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b000001, 
6'b111101, 
6'b111111, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111110, 
6'b000001, 
6'b111110, 
6'b000001, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b111101, 
6'b000001, 
6'b000001, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111110, 
6'b111101, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111101, 
6'b111110, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111101, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111110, 
6'b111110, 
6'b000010, 
6'b111101, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111101, 
6'b111111, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b111101, 
6'b111110, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b000001, 
6'b111101, 
6'b000000, 
6'b000000, 
6'b000010, 
6'b111101, 
6'b111111, 
6'b111101, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b111110, 
6'b000001, 
6'b111111, 
6'b111101, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b000001, 
6'b000001, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b000001, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b111110, 
6'b111110, 
6'b111101, 
6'b111111, 
6'b111111, 
6'b111101, 
6'b000001, 
6'b111110, 
6'b000000, 
6'b111110, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b111110, 
6'b000001, 
6'b000000, 
6'b111111, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b000001, 
6'b000001, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b111101, 
6'b000001, 
6'b000000, 
6'b000001, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b111110, 
6'b111110, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b000001, 
6'b111110, 
6'b111110, 
6'b000001, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b111111, 
6'b111110, 
6'b000001, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111110, 
6'b000010, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111101, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b000001, 
6'b111101, 
6'b111111, 
6'b000001, 
6'b000001, 
6'b111101, 
6'b111110, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b000010, 
6'b000000, 
6'b111101, 
6'b000000, 
6'b111110, 
6'b111110, 
6'b111101, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b111101, 
6'b000000, 
6'b000000, 
6'b111101, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b000001, 
6'b000000, 
6'b111101, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b000010, 
6'b000000, 
6'b000001, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b111101, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111101, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b111110, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b111101, 
6'b111101, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b000001, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b000001, 
6'b000001, 
6'b111110, 
6'b000000, 
6'b000001, 
6'b000001, 
6'b000001, 
6'b111111, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b111110, 
6'b111110, 
6'b000001, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b111101, 
6'b111110, 
6'b111110, 
6'b111111, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111101, 
6'b111111, 
6'b000001, 
6'b000001, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b111101, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111110, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b111110, 
6'b000001, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b111110, 
6'b000001, 
6'b000000, 
6'b111111, 
6'b111110, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b000001, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b000010, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b000010, 
6'b000001, 
6'b111111, 
6'b111101, 
6'b000000, 
6'b111110, 
6'b000010, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111101, 
6'b000000, 
6'b111101, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b111101, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111101, 
6'b111111, 
6'b000001, 
6'b111110, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b111110, 
6'b111111, 
6'b000001, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b111101, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111110, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b111110, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b111101, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b111101, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b111101, 
6'b111101, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111101, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b111101, 
6'b000001, 
6'b111101, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b111110, 
6'b111110, 
6'b111111, 
6'b111101, 
6'b111111, 
6'b111111, 
6'b111110, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b111101, 
6'b000010, 
6'b111111, 
6'b111110, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b111110, 
6'b000001, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b000001, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000010, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b000001, 
6'b111110, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b000010, 
6'b111110, 
6'b000000, 
6'b000001, 
6'b111110, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b111111, 
6'b111110, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111101, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000010, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000001, 
6'b111101, 
6'b000001, 
6'b111111, 
6'b111101, 
6'b111110, 
6'b000010, 
6'b111110, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b000001, 
6'b000001, 
6'b111110, 
6'b000000, 
6'b111101, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b111110, 
6'b000001, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b111101, 
6'b000001, 
6'b111110, 
6'b000001, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b000001, 
6'b111110, 
6'b111110, 
6'b000001, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b000001, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b111101, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b111100, 
6'b111110, 
6'b111110, 
6'b000000, 
6'b111101, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b000001, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b000010, 
6'b111110, 
6'b111110, 
6'b000000, 
6'b000001, 
6'b000001, 
6'b000001, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b000000, 
6'b111110, 
6'b111110, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b111111, 
6'b111101, 
6'b111110, 
6'b000001, 
6'b111110, 
6'b000001, 
6'b000010, 
6'b000001, 
6'b111111, 
6'b111110, 
6'b000000, 
6'b111110, 
6'b111111, 
6'b000000, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000001
};
localparam logic signed [5:0] dlBiases [9:0] = {
6'b000001, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b111111, 
6'b000000, 
6'b111110, 
6'b111111
};
localparam logic signed [5:0] convWeights [0:17] = {
6'b000000, 
6'b000011, 
6'b111110, 
6'b000000, 
6'b000000, 
6'b000100, 
6'b000011, 
6'b000001, 
6'b111110, 
6'b000010, 
6'b111111, 
6'b000001, 
6'b000011, 
6'b000001, 
6'b000011, 
6'b111111, 
6'b000001, 
6'b000000
};
localparam logic signed [5:0] convBiases [1:0] = {
6'b000000, 
6'b000000 
};
endpackage