package data16_8;
localparam logic signed [15:0] dlWeights [0:1279] = {
16'b0000000001000001, 
16'b0000000000000010, 
16'b1111111111001110, 
16'b0000000000000001, 
16'b1111111111101111, 
16'b0000000000100010, 
16'b0000000000010000, 
16'b1111111111001101, 
16'b0000000000001011, 
16'b0000000000101010, 
16'b0000000000101011, 
16'b1111111110111101, 
16'b1111111110011110, 
16'b1111111111010100, 
16'b0000000000011000, 
16'b1111111111100001, 
16'b1111111111101100, 
16'b1111111111111000, 
16'b1111111111110011, 
16'b1111111111111111, 
16'b0000000000011110, 
16'b1111111111000010, 
16'b0000000000001101, 
16'b0000000000010100, 
16'b1111111111110111, 
16'b0000000000000001, 
16'b1111111111101111, 
16'b0000000000001000, 
16'b0000000000010000, 
16'b0000000001000000, 
16'b0000000010010010, 
16'b1111111110010010, 
16'b1111111111000001, 
16'b1111111110110101, 
16'b1111111111000100, 
16'b0000000000011111, 
16'b1111111111111001, 
16'b0000000000101001, 
16'b1111111111101101, 
16'b0000000000110100, 
16'b0000000000100111, 
16'b1111111111011101, 
16'b1111111111111011, 
16'b1111111111010100, 
16'b0000000000000001, 
16'b1111111111100111, 
16'b0000000000101100, 
16'b1111111111011001, 
16'b1111111111100011, 
16'b0000000000000010, 
16'b0000000001011101, 
16'b1111111111011011, 
16'b1111111110111110, 
16'b1111111110101010, 
16'b1111111111010110, 
16'b0000000000011000, 
16'b1111111111111010, 
16'b0000000000100000, 
16'b0000000000010000, 
16'b0000000000011010, 
16'b0000000000111110, 
16'b1111111111001101, 
16'b0000000000010000, 
16'b0000000000010001, 
16'b1111111111010100, 
16'b0000000000111010, 
16'b0000000000110110, 
16'b0000000000000000, 
16'b0000000000101100, 
16'b1111111111101011, 
16'b0000000000000000, 
16'b0000000000110101, 
16'b1111111111000111, 
16'b1111111111011000, 
16'b1111111111010111, 
16'b0000000000011001, 
16'b1111111111110101, 
16'b0000000000101101, 
16'b1111111111000100, 
16'b1111111111010001, 
16'b1111111111101100, 
16'b1111111111100101, 
16'b1111111111000110, 
16'b0000000000011010, 
16'b1111111111011101, 
16'b0000000000100010, 
16'b0000000000000000, 
16'b1111111111010100, 
16'b1111111111110001, 
16'b1111111111100011, 
16'b0000000000001001, 
16'b0000000000000100, 
16'b1111111111100100, 
16'b0000000000000111, 
16'b1111111110111000, 
16'b1111111111110010, 
16'b1111111111000010, 
16'b0000000001010000, 
16'b1111111110111101, 
16'b1111111110110010, 
16'b0000000000000101, 
16'b0000000001001100, 
16'b0000000000000001, 
16'b0000000000001000, 
16'b1111111111011001, 
16'b1111111111111001, 
16'b1111111111010010, 
16'b1111111111010101, 
16'b0000000000011011, 
16'b1111111111001110, 
16'b0000000000000111, 
16'b0000000000101010, 
16'b0000000000001000, 
16'b0000000000100000, 
16'b1111111111000000, 
16'b1111111111100110, 
16'b1111111110111100, 
16'b0000000000011100, 
16'b1111111111010101, 
16'b0000000000010000, 
16'b1111111111010000, 
16'b1111111111110001, 
16'b0000000000000100, 
16'b0000000000010011, 
16'b1111111111000011, 
16'b1111111111101111, 
16'b1111111111000100, 
16'b1111111111100110, 
16'b0000000000000000, 
16'b0000000000010101, 
16'b1111111111010110, 
16'b1111111111101111, 
16'b1111111111100101, 
16'b0000000001000111, 
16'b1111111111010011, 
16'b1111111110101110, 
16'b1111111111011010, 
16'b0000000001010001, 
16'b1111111111110010, 
16'b0000000000001100, 
16'b1111111111111100, 
16'b1111111111101011, 
16'b0000000000000011, 
16'b0000000000001100, 
16'b0000000000110011, 
16'b1111111111110101, 
16'b1111111110111100, 
16'b0000000000110100, 
16'b1111111111110010, 
16'b0000000000010001, 
16'b0000000000000101, 
16'b0000000000010101, 
16'b0000000000100101, 
16'b1111111111111101, 
16'b0000000000010100, 
16'b1111111111011010, 
16'b1111111100111111, 
16'b0000000000110011, 
16'b1111111111110100, 
16'b0000000000011001, 
16'b0000000000101000, 
16'b1111111111110001, 
16'b1111111110111101, 
16'b0000000000101111, 
16'b0000000000110111, 
16'b1111111111100100, 
16'b0000000001000000, 
16'b1111111111110001, 
16'b0000000000001010, 
16'b1111111111111011, 
16'b0000000000100101, 
16'b1111111111111100, 
16'b1111111111110001, 
16'b1111111110101000, 
16'b0000000000000100, 
16'b0000000000001110, 
16'b1111111111101010, 
16'b1111111111111001, 
16'b1111111111100011, 
16'b0000000000100101, 
16'b0000000000111100, 
16'b1111111111000100, 
16'b1111111111111011, 
16'b1111111111101000, 
16'b0000000000111100, 
16'b1111111111111101, 
16'b0000000000100011, 
16'b1111111111100011, 
16'b0000000000110010, 
16'b0000000000000001, 
16'b0000000000111100, 
16'b1111111110100111, 
16'b1111111111011010, 
16'b1111111110111100, 
16'b1111111111111110, 
16'b0000000000010111, 
16'b0000000000001010, 
16'b0000000000011010, 
16'b0000000000100111, 
16'b1111111111110100, 
16'b0000000000110100, 
16'b1111111110111101, 
16'b1111111111100100, 
16'b1111111111011101, 
16'b1111111111111111, 
16'b0000000000000010, 
16'b0000000000000000, 
16'b1111111111110111, 
16'b0000000000000101, 
16'b1111111111100110, 
16'b1111111111110001, 
16'b1111111111110101, 
16'b1111111111110100, 
16'b1111111111001011, 
16'b1111111111111100, 
16'b0000000000000110, 
16'b0000000000110101, 
16'b1111111111101000, 
16'b0000000000000011, 
16'b0000000000001011, 
16'b1111111111011101, 
16'b1111111111110011, 
16'b1111111111001110, 
16'b0000000000101111, 
16'b1111111111001101, 
16'b0000000000111101, 
16'b1111111111010010, 
16'b0000000000000100, 
16'b1111111111101010, 
16'b1111111110111011, 
16'b0000000000101000, 
16'b0000000000111010, 
16'b1111111111001111, 
16'b0000000000010001, 
16'b1111111111111010, 
16'b0000000000000011, 
16'b1111111111100101, 
16'b0000000000101000, 
16'b0000000000001111, 
16'b0000000000001100, 
16'b0000000000000000, 
16'b1111111111100101, 
16'b0000000000010101, 
16'b0000000000011110, 
16'b0000000000010100, 
16'b1111111111101011, 
16'b1111111111010101, 
16'b1111111111101111, 
16'b0000000000011110, 
16'b1111111111011010, 
16'b0000000000010011, 
16'b0000000000010001, 
16'b1111111111101100, 
16'b1111111111011111, 
16'b1111111110111101, 
16'b1111111111100101, 
16'b0000000000000010, 
16'b0000000000000000, 
16'b1111111110110010, 
16'b1111111111001011, 
16'b1111111111000000, 
16'b0000000000001011, 
16'b0000000000000111, 
16'b0000000000010110, 
16'b1111111110101010, 
16'b0000000000000101, 
16'b0000000000011100, 
16'b1111111111001011, 
16'b0000000000000010, 
16'b1111111111111001, 
16'b0000000000000111, 
16'b0000000000101111, 
16'b0000000000001101, 
16'b0000000000000111, 
16'b1111111111110111, 
16'b1111111111001100, 
16'b1111111111000111, 
16'b0000000001000011, 
16'b1111111110111001, 
16'b0000000000000101, 
16'b1111111111111101, 
16'b0000000000000010, 
16'b0000000000010110, 
16'b1111111111110010, 
16'b0000000000001000, 
16'b1111111111100100, 
16'b0000000000011010, 
16'b1111111111111111, 
16'b0000000000100100, 
16'b0000000000010111, 
16'b1111111111100100, 
16'b0000000000011101, 
16'b0000000000011101, 
16'b0000000000000001, 
16'b0000000000010110, 
16'b1111111111100111, 
16'b1111111110110010, 
16'b1111111111111011, 
16'b1111111111010100, 
16'b1111111111101110, 
16'b0000000000001001, 
16'b0000000000110011, 
16'b0000000000001100, 
16'b0000000000010111, 
16'b1111111111101110, 
16'b0000000000001010, 
16'b0000000000010101, 
16'b1111111111101111, 
16'b0000000000011001, 
16'b0000000000110011, 
16'b0000000000011111, 
16'b0000000000010011, 
16'b1111111111110110, 
16'b0000000000001100, 
16'b0000000000100101, 
16'b0000000000010101, 
16'b1111111111000011, 
16'b0000000000000100, 
16'b1111111111110101, 
16'b1111111111111110, 
16'b0000000000100001, 
16'b1111111110111011, 
16'b1111111111011100, 
16'b0000000000011011, 
16'b0000000000110111, 
16'b0000000000000100, 
16'b0000000000110111, 
16'b1111111110111110, 
16'b0000000000000010, 
16'b0000000000011110, 
16'b0000000001000111, 
16'b1111111110111100, 
16'b1111111111101010, 
16'b1111111110101110, 
16'b1111111111110000, 
16'b0000000000011001, 
16'b1111111111011111, 
16'b0000000000001011, 
16'b1111111111101001, 
16'b1111111111011010, 
16'b0000000000011110, 
16'b1111111111101010, 
16'b1111111111110011, 
16'b1111111111010000, 
16'b0000000000001001, 
16'b1111111111101110, 
16'b0000000000001111, 
16'b1111111111100101, 
16'b0000000000101000, 
16'b1111111111011100, 
16'b0000000000101000, 
16'b1111111111101101, 
16'b1111111110100110, 
16'b0000000000001100, 
16'b0000000000100110, 
16'b0000000000000010, 
16'b0000000000000110, 
16'b0000000000001000, 
16'b0000000000101001, 
16'b1111111111100111, 
16'b0000000000001011, 
16'b1111111111000001, 
16'b0000000000100000, 
16'b0000000000100100, 
16'b0000000000000100, 
16'b1111111111101111, 
16'b0000000000010100, 
16'b1111111111110000, 
16'b0000000000010001, 
16'b0000000000001000, 
16'b0000000000000000, 
16'b0000000000000110, 
16'b1111111111011001, 
16'b0000000000001100, 
16'b1111111111110100, 
16'b0000000000001001, 
16'b0000000000110101, 
16'b0000000000100010, 
16'b1111111111111010, 
16'b1111111111001101, 
16'b0000000000011100, 
16'b1111111111000101, 
16'b1111111111101111, 
16'b1111111111100111, 
16'b1111111111111110, 
16'b0000000000101011, 
16'b1111111111110010, 
16'b0000000000000000, 
16'b0000000000111110, 
16'b1111111111110100, 
16'b1111111111110100, 
16'b1111111111101111, 
16'b1111111111111011, 
16'b0000000000100001, 
16'b1111111111010010, 
16'b1111111111101001, 
16'b1111111111101010, 
16'b1111111111001110, 
16'b1111111111011110, 
16'b1111111110111101, 
16'b1111111111100101, 
16'b1111111111100111, 
16'b1111111110111111, 
16'b0000000000110001, 
16'b1111111111001111, 
16'b0000000000010001, 
16'b1111111111010101, 
16'b1111111111010110, 
16'b0000000000011110, 
16'b0000000000000000, 
16'b1111111111010010, 
16'b0000000000001011, 
16'b1111111111001011, 
16'b0000000000101001, 
16'b0000000000010010, 
16'b1111111111101101, 
16'b1111111111011110, 
16'b1111111111100000, 
16'b0000000000011001, 
16'b1111111111010000, 
16'b0000000000000010, 
16'b0000000000101001, 
16'b0000000000010110, 
16'b0000000000011011, 
16'b1111111111010011, 
16'b0000000000110011, 
16'b0000000000100111, 
16'b0000000000000110, 
16'b0000000000111010, 
16'b0000000000000111, 
16'b1111111110111001, 
16'b0000000000110110, 
16'b0000000000010100, 
16'b0000000000101100, 
16'b1111111111000111, 
16'b1111111111110100, 
16'b0000000000001110, 
16'b1111111111010011, 
16'b1111111111011001, 
16'b1111111111011011, 
16'b1111111111100101, 
16'b0000000000111010, 
16'b0000000000000011, 
16'b0000000000011010, 
16'b0000000000000011, 
16'b0000000000110000, 
16'b0000000000101110, 
16'b1111111111000011, 
16'b1111111111010110, 
16'b0000000000100011, 
16'b1111111111011110, 
16'b1111111111110110, 
16'b1111111111110110, 
16'b0000000000100000, 
16'b0000000000001100, 
16'b1111111111111101, 
16'b1111111111010101, 
16'b0000000000100111, 
16'b1111111111110010, 
16'b0000000000101011, 
16'b0000000000001111, 
16'b0000000000010101, 
16'b1111111111101111, 
16'b0000000000000100, 
16'b0000000000101011, 
16'b1111111111110111, 
16'b1111111111111101, 
16'b1111111111111010, 
16'b1111111111011001, 
16'b0000000001000000, 
16'b0000000000001001, 
16'b1111111111100001, 
16'b1111111111111010, 
16'b0000000000001110, 
16'b1111111111110100, 
16'b1111111111110100, 
16'b0000000000001001, 
16'b0000000000110010, 
16'b0000000000011100, 
16'b0000000000101101, 
16'b0000000000001111, 
16'b1111111111011010, 
16'b0000000000001010, 
16'b1111111111011010, 
16'b1111111111101010, 
16'b1111111111100001, 
16'b0000000000000000, 
16'b0000000000000101, 
16'b0000000000010101, 
16'b0000000000001100, 
16'b0000000000010000, 
16'b1111111110110011, 
16'b1111111111011000, 
16'b1111111111111000, 
16'b0000000000000111, 
16'b0000000000111101, 
16'b0000000000111100, 
16'b1111111110111100, 
16'b1111111111110111, 
16'b0000000000100001, 
16'b0000000000110101, 
16'b1111111110111100, 
16'b1111111111011010, 
16'b0000000000000111, 
16'b0000000000100101, 
16'b1111111111101000, 
16'b1111111111101110, 
16'b1111111111110010, 
16'b1111111111111101, 
16'b0000000000110101, 
16'b0000000000101010, 
16'b1111111111111011, 
16'b1111111111101101, 
16'b0000000000100101, 
16'b0000000000010010, 
16'b0000000000100010, 
16'b1111111111111001, 
16'b1111111111100001, 
16'b1111111111110001, 
16'b1111111111111001, 
16'b1111111111001010, 
16'b0000000000001011, 
16'b1111111111001100, 
16'b0000000000011001, 
16'b1111111111111000, 
16'b1111111111111001, 
16'b0000000000100000, 
16'b0000000000000100, 
16'b1111111111111010, 
16'b0000000000010101, 
16'b0000000000010000, 
16'b0000000000001101, 
16'b0000000000000110, 
16'b0000000000011000, 
16'b1111111111011111, 
16'b0000000001000000, 
16'b0000000000011111, 
16'b1111111110111010, 
16'b0000000000000100, 
16'b1111111111001000, 
16'b1111111111000110, 
16'b1111111110110101, 
16'b1111111111110010, 
16'b1111111111101010, 
16'b1111111111100000, 
16'b0000000000010110, 
16'b0000000000000100, 
16'b1111111111001111, 
16'b0000000000001010, 
16'b1111111111100001, 
16'b1111111111100100, 
16'b1111111111101000, 
16'b1111111111101111, 
16'b1111111111100110, 
16'b0000000000000100, 
16'b1111111111110010, 
16'b0000000000100101, 
16'b1111111111100000, 
16'b0000000000001101, 
16'b0000000000000110, 
16'b0000000000010110, 
16'b0000000000110110, 
16'b0000000000000000, 
16'b1111111111011101, 
16'b1111111111101000, 
16'b0000000000011100, 
16'b0000000000100011, 
16'b1111111110101111, 
16'b0000000000010011, 
16'b0000000000000100, 
16'b1111111110111010, 
16'b0000000000101101, 
16'b1111111111101100, 
16'b0000000000000001, 
16'b1111111111011011, 
16'b0000000000101100, 
16'b0000000000011111, 
16'b1111111110100110, 
16'b0000000000100011, 
16'b0000000000010111, 
16'b0000000000010110, 
16'b0000000001001010, 
16'b0000000000010100, 
16'b0000000000101000, 
16'b1111111111011000, 
16'b0000000000001001, 
16'b1111111111110001, 
16'b0000000000010001, 
16'b0000000000111011, 
16'b0000000000011101, 
16'b1111111110101110, 
16'b0000000000101001, 
16'b1111111111101101, 
16'b0000000000001011, 
16'b1111111111011111, 
16'b1111111111010010, 
16'b0000000000001000, 
16'b0000000000011110, 
16'b0000000000001111, 
16'b1111111111110001, 
16'b1111111110110110, 
16'b0000000000010010, 
16'b0000000000000110, 
16'b0000000000100101, 
16'b0000000000000001, 
16'b0000000000001000, 
16'b0000000000100111, 
16'b0000000000100010, 
16'b1111111111101101, 
16'b0000000000011011, 
16'b1111111111011111, 
16'b1111111111011111, 
16'b1111111111101010, 
16'b0000000000101100, 
16'b1111111111100001, 
16'b1111111111010011, 
16'b0000000000000111, 
16'b0000000000011011, 
16'b0000000000100010, 
16'b1111111111100111, 
16'b1111111110111011, 
16'b1111111110111001, 
16'b0000000000011110, 
16'b0000000000000011, 
16'b0000000000101011, 
16'b0000000000100011, 
16'b0000000000011101, 
16'b0000000000101110, 
16'b1111111111101001, 
16'b1111111111111100, 
16'b0000000000001011, 
16'b0000000000010010, 
16'b0000000000100111, 
16'b0000000000101011, 
16'b0000000000110100, 
16'b1111111111011110, 
16'b0000000000000000, 
16'b0000000000110101, 
16'b0000000000100110, 
16'b0000000000100100, 
16'b1111111111111100, 
16'b1111111111010111, 
16'b1111111111110101, 
16'b1111111111110110, 
16'b1111111111011110, 
16'b1111111111000001, 
16'b0000000000100001, 
16'b0000000000011110, 
16'b0000000000101000, 
16'b0000000000000000, 
16'b1111111111100111, 
16'b1111111111110101, 
16'b1111111111100001, 
16'b0000000000000111, 
16'b0000000000000000, 
16'b0000000000101111, 
16'b0000000000010100, 
16'b1111111110111000, 
16'b1111111111011011, 
16'b1111111111010010, 
16'b1111111111111110, 
16'b1111111111000110, 
16'b1111111111110011, 
16'b1111111111101101, 
16'b0000000000001101, 
16'b0000000000000010, 
16'b0000000000001000, 
16'b1111111110110011, 
16'b1111111111111101, 
16'b0000000000100010, 
16'b0000000000110110, 
16'b1111111111111010, 
16'b1111111111000011, 
16'b0000000000011110, 
16'b1111111111110001, 
16'b0000000000101101, 
16'b1111111111111110, 
16'b1111111110110111, 
16'b1111111111101000, 
16'b0000000000000101, 
16'b1111111111000100, 
16'b1111111111111010, 
16'b0000000000101101, 
16'b1111111111101101, 
16'b1111111111111101, 
16'b0000000000101011, 
16'b0000000000001110, 
16'b1111111111101101, 
16'b0000000000101110, 
16'b1111111111101110, 
16'b0000000000010011, 
16'b0000000000000011, 
16'b1111111111001110, 
16'b0000000000101000, 
16'b1111111111100110, 
16'b0000000000000010, 
16'b0000000000000101, 
16'b1111111111101001, 
16'b1111111111110011, 
16'b0000000000011100, 
16'b0000000000000000, 
16'b0000000000001011, 
16'b0000000000010011, 
16'b1111111111100011, 
16'b0000000000001110, 
16'b1111111111010101, 
16'b1111111111111110, 
16'b1111111111100110, 
16'b1111111111100101, 
16'b1111111111011001, 
16'b0000000000000110, 
16'b0000000000010101, 
16'b0000000000001011, 
16'b1111111111101100, 
16'b1111111111011010, 
16'b0000000000101010, 
16'b1111111111100111, 
16'b0000000000000000, 
16'b0000000000110011, 
16'b0000000000000001, 
16'b1111111111001100, 
16'b0000000000100011, 
16'b1111111111011100, 
16'b0000000000010111, 
16'b0000000000001111, 
16'b0000000000010000, 
16'b0000000000100001, 
16'b1111111111011000, 
16'b0000000000001100, 
16'b1111111111100110, 
16'b1111111111010001, 
16'b0000000000011011, 
16'b1111111111001110, 
16'b0000000000101101, 
16'b0000000000001000, 
16'b1111111111101110, 
16'b1111111111001100, 
16'b1111111111101001, 
16'b0000000000101010, 
16'b1111111111100000, 
16'b0000000000000010, 
16'b1111111111101010, 
16'b0000000000110000, 
16'b1111111111110111, 
16'b0000000000000100, 
16'b0000000000011000, 
16'b1111111111100110, 
16'b1111111111100011, 
16'b0000000000001100, 
16'b0000000000000110, 
16'b1111111111000101, 
16'b0000000000110110, 
16'b1111111111110100, 
16'b0000000000110010, 
16'b0000000000011100, 
16'b0000000000011001, 
16'b1111111111011100, 
16'b1111111111110100, 
16'b1111111111110100, 
16'b1111111111101110, 
16'b1111111111111010, 
16'b0000000000011100, 
16'b1111111111100000, 
16'b0000000000011001, 
16'b0000000000000101, 
16'b0000000000001000, 
16'b0000000000011010, 
16'b0000000000101000, 
16'b0000000000010101, 
16'b1111111111100010, 
16'b0000000000001110, 
16'b1111111111000011, 
16'b0000000000010001, 
16'b1111111111101101, 
16'b0000000000011000, 
16'b1111111111101001, 
16'b1111111111100100, 
16'b0000000000010101, 
16'b1111111111011000, 
16'b1111111111100111, 
16'b1111111111010100, 
16'b0000000000000111, 
16'b1111111111100011, 
16'b0000000000111001, 
16'b1111111111111010, 
16'b1111111111100010, 
16'b1111111111111111, 
16'b0000000000010100, 
16'b0000000000010100, 
16'b0000000000101011, 
16'b1111111111101011, 
16'b1111111111010000, 
16'b0000000000000011, 
16'b1111111111011110, 
16'b1111111111101011, 
16'b1111111111001000, 
16'b0000000000011011, 
16'b0000000001000011, 
16'b0000000000011001, 
16'b0000000000101001, 
16'b1111111111111110, 
16'b1111111111100011, 
16'b0000000000100100, 
16'b1111111111110000, 
16'b0000000000101000, 
16'b1111111111101100, 
16'b0000000000001011, 
16'b1111111111010001, 
16'b0000000001000110, 
16'b0000000000111100, 
16'b1111111111100100, 
16'b1111111110101110, 
16'b0000000000000101, 
16'b1111111111011000, 
16'b0000000001000000, 
16'b1111111111111000, 
16'b1111111111100110, 
16'b0000000000000110, 
16'b1111111111100011, 
16'b1111111111100101, 
16'b1111111111101110, 
16'b1111111110110011, 
16'b0000000000000111, 
16'b1111111110110101, 
16'b1111111111101010, 
16'b0000000000000110, 
16'b0000000000010111, 
16'b1111111111100011, 
16'b1111111111111011, 
16'b0000000000001010, 
16'b1111111111101101, 
16'b1111111110101010, 
16'b1111111111101101, 
16'b0000000000001101, 
16'b0000000000001001, 
16'b0000000000010010, 
16'b0000000000010100, 
16'b1111111110111011, 
16'b1111111111101000, 
16'b0000000000101100, 
16'b1111111111001110, 
16'b1111111111101110, 
16'b0000000000111011, 
16'b1111111111100110, 
16'b0000000000000001, 
16'b1111111111100111, 
16'b0000000000001000, 
16'b1111111111110101, 
16'b1111111111101110, 
16'b0000000000101111, 
16'b1111111111001111, 
16'b1111111111101110, 
16'b0000000000100100, 
16'b0000000000101110, 
16'b1111111111110010, 
16'b0000000000010000, 
16'b1111111111110110, 
16'b1111111110111010, 
16'b1111111111101111, 
16'b0000000000001001, 
16'b1111111111100111, 
16'b1111111111111110, 
16'b1111111111110000, 
16'b1111111111100111, 
16'b0000000000100110, 
16'b1111111111100111, 
16'b1111111111100000, 
16'b0000000000000011, 
16'b1111111111110000, 
16'b0000000000010100, 
16'b1111111111010110, 
16'b0000000000101000, 
16'b0000000000011111, 
16'b0000000000000010, 
16'b1111111111111110, 
16'b1111111111011100, 
16'b1111111111010101, 
16'b1111111111100011, 
16'b1111111111101101, 
16'b1111111111110111, 
16'b0000000000001010, 
16'b0000000000111100, 
16'b1111111111101110, 
16'b1111111111000111, 
16'b0000000000111010, 
16'b1111111111100011, 
16'b1111111111111001, 
16'b0000000000001000, 
16'b0000000000011010, 
16'b1111111111011111, 
16'b1111111111100010, 
16'b1111111111110011, 
16'b0000000000011101, 
16'b1111111111100111, 
16'b0000000000011001, 
16'b0000000000011101, 
16'b1111111111010011, 
16'b0000000000000001, 
16'b0000000000000000, 
16'b1111111111110011, 
16'b1111111111101100, 
16'b0000000000000101, 
16'b1111111111110011, 
16'b0000000000001110, 
16'b0000000000001101, 
16'b1111111111010100, 
16'b1111111111100010, 
16'b0000000000000111, 
16'b0000000000011110, 
16'b1111111111001000, 
16'b1111111110111001, 
16'b1111111111100111, 
16'b1111111111110100, 
16'b1111111111110111, 
16'b1111111111111011, 
16'b1111111111011011, 
16'b0000000000010101, 
16'b0000000000010111, 
16'b1111111111100111, 
16'b0000000000011011, 
16'b1111111111111100, 
16'b1111111111101110, 
16'b0000000000101100, 
16'b1111111111100001, 
16'b1111111111110110, 
16'b1111111111100001, 
16'b0000000000001100, 
16'b0000000000100100, 
16'b1111111111111110, 
16'b0000000000010110, 
16'b1111111110110111, 
16'b0000000000000110, 
16'b1111111111100101, 
16'b1111111111101011, 
16'b0000000000100110, 
16'b1111111111010001, 
16'b0000000000010101, 
16'b1111111111101011, 
16'b0000000000000001, 
16'b0000000000000001, 
16'b1111111111001100, 
16'b1111111111111100, 
16'b0000000000000111, 
16'b1111111111011011, 
16'b0000000000001000, 
16'b0000000000101000, 
16'b1111111111100100, 
16'b0000000000011110, 
16'b1111111111110001, 
16'b0000000000110111, 
16'b1111111110101111, 
16'b1111111110101100, 
16'b0000000000011000, 
16'b1111111111101001, 
16'b0000000000001010, 
16'b1111111111011101, 
16'b1111111111110101, 
16'b0000000000011101, 
16'b0000000000001000, 
16'b1111111111111110, 
16'b0000000000001000, 
16'b1111111111100100, 
16'b0000000000100010, 
16'b1111111111111110, 
16'b1111111111100111, 
16'b0000000000010100, 
16'b1111111111111000, 
16'b0000000000000011, 
16'b0000000000011111, 
16'b1111111111001001, 
16'b1111111111100000, 
16'b1111111110101111, 
16'b0000000000010000, 
16'b1111111111001001, 
16'b0000000000011000, 
16'b0000000000010011, 
16'b1111111111111111, 
16'b1111111111011111, 
16'b1111111111100101, 
16'b0000000000011100, 
16'b1111111111111010, 
16'b1111111110111111, 
16'b0000000000110010, 
16'b1111111110111000, 
16'b1111111111011001, 
16'b1111111111111000, 
16'b0000000000000000, 
16'b1111111111010010, 
16'b1111111111101011, 
16'b1111111111111111, 
16'b1111111111111011, 
16'b1111111111110100, 
16'b1111111111111101, 
16'b1111111111100010, 
16'b0000000000111000, 
16'b1111111111110001, 
16'b0000000000000111, 
16'b0000000000000111, 
16'b1111111111110110, 
16'b0000000000001010, 
16'b0000000000000101, 
16'b1111111111110011, 
16'b1111111111110100, 
16'b0000000000001101, 
16'b0000000000000110, 
16'b0000000000001011, 
16'b0000000000010101, 
16'b1111111111011010, 
16'b0000000000111110, 
16'b1111111111101000, 
16'b0000000000001000, 
16'b1111111111101010, 
16'b0000000000010100, 
16'b1111111111010011, 
16'b1111111111011100, 
16'b1111111111000111, 
16'b1111111111110101, 
16'b1111111110101100, 
16'b1111111111111101, 
16'b1111111111100011, 
16'b1111111111010010, 
16'b1111111111011110, 
16'b1111111111101111, 
16'b1111111111100010, 
16'b0000000000101010, 
16'b1111111110101111, 
16'b0000000001000010, 
16'b1111111111110101, 
16'b1111111111011110, 
16'b1111111111110101, 
16'b1111111111001110, 
16'b0000000000001001, 
16'b0000000000010110, 
16'b1111111111010101, 
16'b0000000000001011, 
16'b1111111111000100, 
16'b0000000000100001, 
16'b1111111111001111, 
16'b0000000000001011, 
16'b1111111111101000, 
16'b1111111111110000, 
16'b0000000000101100, 
16'b0000000000100100, 
16'b1111111111100110, 
16'b0000000000100011, 
16'b0000000000001110, 
16'b0000000000001001, 
16'b0000000000110110, 
16'b0000000000011111, 
16'b1111111111100100, 
16'b1111111111100000, 
16'b0000000000101110, 
16'b0000000000101010, 
16'b0000000000000011, 
16'b0000000000011000, 
16'b0000000000001011, 
16'b0000000000001011, 
16'b1111111111110110, 
16'b0000000000100111, 
16'b1111111111111000, 
16'b0000000000000000, 
16'b0000000000001111, 
16'b0000000001001100, 
16'b1111111111010101, 
16'b1111111111101110, 
16'b0000000000000001, 
16'b0000000000100000, 
16'b0000000000100111, 
16'b1111111111011000, 
16'b1111111111010110, 
16'b0000000000000101, 
16'b0000000000001110, 
16'b0000000000000101, 
16'b0000000000001000, 
16'b0000000000010010, 
16'b0000000000001110, 
16'b0000000000100001, 
16'b1111111111111110, 
16'b0000000000000101, 
16'b0000000000100100, 
16'b1111111111111101, 
16'b1111111111110100, 
16'b0000000000001000, 
16'b1111111111001100, 
16'b0000000000000110, 
16'b0000000000010110, 
16'b1111111111010111, 
16'b0000000000111110, 
16'b1111111111111100, 
16'b0000000000001111, 
16'b1111111111111101, 
16'b1111111111110110, 
16'b1111111111110100, 
16'b0000000000011101, 
16'b0000000000111111, 
16'b0000000000000000, 
16'b0000000000011000, 
16'b0000000001000000, 
16'b1111111111001111, 
16'b0000000000011110, 
16'b0000000000100000, 
16'b1111111111011110, 
16'b0000000000000111, 
16'b0000000000100111, 
16'b0000000000000011, 
16'b0000000000011101, 
16'b1111111111111011, 
16'b0000000000110111, 
16'b0000000000010111, 
16'b1111111111101000, 
16'b1111111111000011, 
16'b1111111111011011, 
16'b0000000000001100, 
16'b0000000000000011, 
16'b1111111111111000, 
16'b0000000000010001, 
16'b0000000000010110, 
16'b0000000000010101, 
16'b1111111111000110, 
16'b0000000000001011, 
16'b0000000000011010, 
16'b1111111111001101, 
16'b1111111111100101, 
16'b1111111111110111, 
16'b0000000000110010, 
16'b0000000000110101, 
16'b1111111111111111, 
16'b0000000000011101, 
16'b1111111111001101, 
16'b1111111111101101, 
16'b1111111111101111, 
16'b1111111111111001, 
16'b0000000000000100, 
16'b1111111110111100, 
16'b0000000000011101, 
16'b1111111111110010, 
16'b1111111111110010, 
16'b1111111111010100, 
16'b0000000000000111, 
16'b1111111111111101, 
16'b0000000001001011, 
16'b1111111111000101, 
16'b0000000000010000, 
16'b0000000000000001, 
16'b1111111111100001, 
16'b1111111111101100, 
16'b0000000000001010, 
16'b1111111111010101, 
16'b1111111111100111, 
16'b1111111111000111, 
16'b1111111111110001, 
16'b0000000000011011, 
16'b0000000000110011, 
16'b1111111111011110, 
16'b1111111111110011, 
16'b0000000000001001, 
16'b0000000000101001, 
16'b1111111111101111, 
16'b1111111111111111, 
16'b1111111111111010, 
16'b0000000000101100, 
16'b1111111110111011, 
16'b0000000000101010, 
16'b1111111111100100, 
16'b1111111110111110, 
16'b1111111111011110, 
16'b0000000001000010, 
16'b1111111111001011, 
16'b1111111111110001, 
16'b1111111111000000, 
16'b0000000000011000, 
16'b0000000000111000, 
16'b0000000000111011, 
16'b1111111111011111, 
16'b0000000000000011, 
16'b1111111110111100, 
16'b0000000000011011, 
16'b1111111111100001, 
16'b0000000000100101, 
16'b0000000000000001, 
16'b0000000000010100, 
16'b1111111111100000, 
16'b1111111111100110, 
16'b1111111111011101, 
16'b0000000000001100, 
16'b0000000000010001, 
16'b0000000000110111, 
16'b0000000000001000, 
16'b1111111111100001, 
16'b1111111111110000, 
16'b1111111111001001, 
16'b0000000000101010, 
16'b0000000000011101, 
16'b1111111111010001, 
16'b1111111111110011, 
16'b1111111110111100, 
16'b0000000000101010, 
16'b1111111111001100, 
16'b0000000000110100, 
16'b1111111111011111, 
16'b0000000000001100, 
16'b0000000000000110, 
16'b0000000000101000, 
16'b1111111111011011, 
16'b1111111111010111, 
16'b0000000000101101, 
16'b1111111111100110, 
16'b0000000000000101, 
16'b1111111111010101, 
16'b0000000000000011, 
16'b1111111111101000, 
16'b0000000000011101, 
16'b1111111111101101, 
16'b1111111111100110, 
16'b1111111111101000, 
16'b0000000000011001, 
16'b1111111111101100, 
16'b1111111111110101, 
16'b0000000000010100, 
16'b0000000000100110, 
16'b1111111111000010, 
16'b0000000000000100, 
16'b0000000000000110, 
16'b1111111110111110, 
16'b1111111111110110, 
16'b0000000000110001, 
16'b0000000000011101, 
16'b1111111111000111, 
16'b0000000000011110, 
16'b1111111110010001, 
16'b1111111111001011, 
16'b1111111111010010, 
16'b0000000000000100, 
16'b1111111110111010, 
16'b1111111111101110, 
16'b0000000000000100, 
16'b1111111111101000, 
16'b0000000000111111, 
16'b0000000000001000, 
16'b0000000000000010, 
16'b0000000000000000, 
16'b0000000001001011, 
16'b1111111111010011, 
16'b1111111111010111, 
16'b0000000000001011, 
16'b0000000000101010, 
16'b0000000000100000, 
16'b0000000000100000, 
16'b1111111111100010, 
16'b1111111111010111, 
16'b0000000000000111, 
16'b1111111111011101, 
16'b0000000000001010, 
16'b0000000000001111, 
16'b0000000000000101, 
16'b1111111111000101, 
16'b1111111111000101, 
16'b1111111111111001, 
16'b1111111111110001, 
16'b1111111111110110, 
16'b1111111111000001, 
16'b0000000000001010, 
16'b1111111111101010, 
16'b1111111110110101, 
16'b1111111111011110, 
16'b0000000000101011, 
16'b1111111111001111, 
16'b0000000000100100, 
16'b0000000001000000, 
16'b0000000000111111, 
16'b1111111111111110, 
16'b1111111111010101, 
16'b0000000000011011, 
16'b1111111111010110, 
16'b1111111111101110, 
16'b0000000000011001, 
16'b1111111111111001, 
16'b1111111111110111, 
16'b1111111111110110, 
16'b0000000000100000

};
localparam logic signed [15:0] dlBiases [9:0] = {
16'b0000000000101010, 
16'b1111111111111111, 
16'b1111111111111111, 
16'b1111111111110001, 
16'b1111111111110000, 
16'b1111111111111010, 
16'b1111111111111010, 
16'b0000000000010011, 
16'b1111111111010001, 
16'b1111111111111010 

};
localparam logic signed [15:0] convWeights [0:17] = {
16'b0000000000011100, 
16'b0000000001111011, 
16'b1111111111000010, 
16'b0000000000010111, 
16'b0000000000000011, 
16'b0000000010000011, 
16'b0000000001100111, 
16'b0000000000110011, 
16'b1111111111000101, 
16'b0000000001011001, 
16'b1111111111101001, 
16'b0000000000110101, 
16'b0000000001111111, 
16'b0000000000101000, 
16'b0000000001100010, 
16'b1111111111111101, 
16'b0000000000101110, 
16'b0000000000011101

};
localparam logic signed [15:0] convBiases [1:0] = {
16'b0000000000000000, 
16'b0000000000000000
};
endpackage