package data20_10;
localparam logic signed [19:0] dlWeights [0:1279] = {
20'b00000000000100000111, 
20'b00000000000000001010, 
20'b11111111111100111000, 
20'b00000000000000000110, 
20'b11111111111110111101, 
20'b00000000000010001001, 
20'b00000000000001000000, 
20'b11111111111100110100, 
20'b00000000000000101110, 
20'b00000000000010101011, 
20'b00000000000010101100, 
20'b11111111111011110111, 
20'b11111111111001111011, 
20'b11111111111101010011, 
20'b00000000000001100010, 
20'b11111111111110000100, 
20'b11111111111110110011, 
20'b11111111111111100001, 
20'b11111111111111001100, 
20'b11111111111111111100, 
20'b00000000000001111011, 
20'b11111111111100001011, 
20'b00000000000000110111, 
20'b00000000000001010010, 
20'b11111111111111011110, 
20'b00000000000000000101, 
20'b11111111111110111100, 
20'b00000000000000100011, 
20'b00000000000001000010, 
20'b00000000000100000011, 
20'b00000000001001001011, 
20'b11111111111001001010, 
20'b11111111111100000110, 
20'b11111111111011010100, 
20'b11111111111100010001, 
20'b00000000000001111100, 
20'b11111111111111100101, 
20'b00000000000010100110, 
20'b11111111111110110111, 
20'b00000000000011010010, 
20'b00000000000010011111, 
20'b11111111111101110101, 
20'b11111111111111101110, 
20'b11111111111101010010, 
20'b00000000000000000101, 
20'b11111111111110011110, 
20'b00000000000010110010, 
20'b11111111111101100110, 
20'b11111111111110001101, 
20'b00000000000000001010, 
20'b00000000000101110101, 
20'b11111111111101101101, 
20'b11111111111011111000, 
20'b11111111111010101001, 
20'b11111111111101011010, 
20'b00000000000001100011, 
20'b11111111111111101001, 
20'b00000000000010000010, 
20'b00000000000001000001, 
20'b00000000000001101001, 
20'b00000000000011111000, 
20'b11111111111100110101, 
20'b00000000000001000011, 
20'b00000000000001000100, 
20'b11111111111101010010, 
20'b00000000000011101001, 
20'b00000000000011011010, 
20'b00000000000000000010, 
20'b00000000000010110011, 
20'b11111111111110101110, 
20'b00000000000000000011, 
20'b00000000000011010110, 
20'b11111111111100011111, 
20'b11111111111101100011, 
20'b11111111111101011101, 
20'b00000000000001100101, 
20'b11111111111111010111, 
20'b00000000000010110100, 
20'b11111111111100010001, 
20'b11111111111101000111, 
20'b11111111111110110010, 
20'b11111111111110010100, 
20'b11111111111100011000, 
20'b00000000000001101011, 
20'b11111111111101110110, 
20'b00000000000010001000, 
20'b00000000000000000000, 
20'b11111111111101010011, 
20'b11111111111111000111, 
20'b11111111111110001110, 
20'b00000000000000100100, 
20'b00000000000000010001, 
20'b11111111111110010011, 
20'b00000000000000011100, 
20'b11111111111011100000, 
20'b11111111111111001011, 
20'b11111111111100001011, 
20'b00000000000101000001, 
20'b11111111111011110110, 
20'b11111111111011001010, 
20'b00000000000000010101, 
20'b00000000000100110000, 
20'b00000000000000000101, 
20'b00000000000000100011, 
20'b11111111111101100110, 
20'b11111111111111100111, 
20'b11111111111101001001, 
20'b11111111111101010100, 
20'b00000000000001101111, 
20'b11111111111100111000, 
20'b00000000000000011100, 
20'b00000000000010101010, 
20'b00000000000000100011, 
20'b00000000000010000010, 
20'b11111111111100000010, 
20'b11111111111110011001, 
20'b11111111111011110010, 
20'b00000000000001110001, 
20'b11111111111101010111, 
20'b00000000000001000001, 
20'b11111111111101000001, 
20'b11111111111111000111, 
20'b00000000000000010001, 
20'b00000000000001001101, 
20'b11111111111100001110, 
20'b11111111111110111101, 
20'b11111111111100010010, 
20'b11111111111110011000, 
20'b00000000000000000010, 
20'b00000000000001010100, 
20'b11111111111101011010, 
20'b11111111111110111110, 
20'b11111111111110010101, 
20'b00000000000100011110, 
20'b11111111111101001101, 
20'b11111111111010111000, 
20'b11111111111101101001, 
20'b00000000000101000100, 
20'b11111111111111001001, 
20'b00000000000000110000, 
20'b11111111111111110011, 
20'b11111111111110101111, 
20'b00000000000000001111, 
20'b00000000000000110000, 
20'b00000000000011001111, 
20'b11111111111111010110, 
20'b11111111111011110010, 
20'b00000000000011010011, 
20'b11111111111111001000, 
20'b00000000000001000110, 
20'b00000000000000010100, 
20'b00000000000001010101, 
20'b00000000000010010101, 
20'b11111111111111110101, 
20'b00000000000001010011, 
20'b11111111111101101010, 
20'b11111111110011111111, 
20'b00000000000011001100, 
20'b11111111111111010010, 
20'b00000000000001100110, 
20'b00000000000010100011, 
20'b11111111111111000100, 
20'b11111111111011110111, 
20'b00000000000010111101, 
20'b00000000000011011100, 
20'b11111111111110010011, 
20'b00000000000100000010, 
20'b11111111111111000101, 
20'b00000000000000101011, 
20'b11111111111111101100, 
20'b00000000000010010111, 
20'b11111111111111110000, 
20'b11111111111111000100, 
20'b11111111111010100010, 
20'b00000000000000010011, 
20'b00000000000000111001, 
20'b11111111111110101011, 
20'b11111111111111100100, 
20'b11111111111110001101, 
20'b00000000000010010110, 
20'b00000000000011110000, 
20'b11111111111100010000, 
20'b11111111111111101110, 
20'b11111111111110100010, 
20'b00000000000011110010, 
20'b11111111111111110110, 
20'b00000000000010001110, 
20'b11111111111110001111, 
20'b00000000000011001011, 
20'b00000000000000000111, 
20'b00000000000011110000, 
20'b11111111111010011100, 
20'b11111111111101101011, 
20'b11111111111011110001, 
20'b11111111111111111001, 
20'b00000000000001011101, 
20'b00000000000000101011, 
20'b00000000000001101010, 
20'b00000000000010011111, 
20'b11111111111111010010, 
20'b00000000000011010001, 
20'b11111111111011110100, 
20'b11111111111110010010, 
20'b11111111111101110100, 
20'b11111111111111111110, 
20'b00000000000000001011, 
20'b00000000000000000011, 
20'b11111111111111011111, 
20'b00000000000000010101, 
20'b11111111111110011000, 
20'b11111111111111000101, 
20'b11111111111111010101, 
20'b11111111111111010010, 
20'b11111111111100101100, 
20'b11111111111111110000, 
20'b00000000000000011010, 
20'b00000000000011010100, 
20'b11111111111110100010, 
20'b00000000000000001111, 
20'b00000000000000101101, 
20'b11111111111101110111, 
20'b11111111111111001100, 
20'b11111111111100111011, 
20'b00000000000010111110, 
20'b11111111111100110111, 
20'b00000000000011110101, 
20'b11111111111101001001, 
20'b00000000000000010011, 
20'b11111111111110101011, 
20'b11111111111011101111, 
20'b00000000000010100010, 
20'b00000000000011101011, 
20'b11111111111100111111, 
20'b00000000000001000111, 
20'b11111111111111101000, 
20'b00000000000000001110, 
20'b11111111111110010100, 
20'b00000000000010100010, 
20'b00000000000000111111, 
20'b00000000000000110011, 
20'b00000000000000000011, 
20'b11111111111110010100, 
20'b00000000000001010100, 
20'b00000000000001111011, 
20'b00000000000001010000, 
20'b11111111111110101100, 
20'b11111111111101010110, 
20'b11111111111110111110, 
20'b00000000000001111001, 
20'b11111111111101101001, 
20'b00000000000001001100, 
20'b00000000000001000110, 
20'b11111111111110110011, 
20'b11111111111101111111, 
20'b11111111111011110100, 
20'b11111111111110010110, 
20'b00000000000000001010, 
20'b00000000000000000001, 
20'b11111111111011001010, 
20'b11111111111100101111, 
20'b11111111111100000000, 
20'b00000000000000101100, 
20'b00000000000000011111, 
20'b00000000000001011010, 
20'b11111111111010101011, 
20'b00000000000000010111, 
20'b00000000000001110001, 
20'b11111111111100101110, 
20'b00000000000000001001, 
20'b11111111111111100111, 
20'b00000000000000011110, 
20'b00000000000010111100, 
20'b00000000000000110100, 
20'b00000000000000011101, 
20'b11111111111111011100, 
20'b11111111111100110001, 
20'b11111111111100011100, 
20'b00000000000100001111, 
20'b11111111111011100101, 
20'b00000000000000010101, 
20'b11111111111111110100, 
20'b00000000000000001000, 
20'b00000000000001011010, 
20'b11111111111111001010, 
20'b00000000000000100011, 
20'b11111111111110010000, 
20'b00000000000001101000, 
20'b11111111111111111110, 
20'b00000000000010010001, 
20'b00000000000001011101, 
20'b11111111111110010001, 
20'b00000000000001110110, 
20'b00000000000001110111, 
20'b00000000000000000101, 
20'b00000000000001011010, 
20'b11111111111110011110, 
20'b11111111111011001000, 
20'b11111111111111101101, 
20'b11111111111101010001, 
20'b11111111111110111010, 
20'b00000000000000100110, 
20'b00000000000011001100, 
20'b00000000000000110000, 
20'b00000000000001011110, 
20'b11111111111110111000, 
20'b00000000000000101000, 
20'b00000000000001010101, 
20'b11111111111110111100, 
20'b00000000000001100110, 
20'b00000000000011001110, 
20'b00000000000001111111, 
20'b00000000000001001100, 
20'b11111111111111011001, 
20'b00000000000000110000, 
20'b00000000000010010111, 
20'b00000000000001010100, 
20'b11111111111100001101, 
20'b00000000000000010010, 
20'b11111111111111010100, 
20'b11111111111111111011, 
20'b00000000000010000101, 
20'b11111111111011101101, 
20'b11111111111101110011, 
20'b00000000000001101100, 
20'b00000000000011011100, 
20'b00000000000000010011, 
20'b00000000000011011111, 
20'b11111111111011111001, 
20'b00000000000000001000, 
20'b00000000000001111010, 
20'b00000000000100011101, 
20'b11111111111011110001, 
20'b11111111111110101000, 
20'b11111111111010111011, 
20'b11111111111111000000, 
20'b00000000000001100111, 
20'b11111111111101111111, 
20'b00000000000000101100, 
20'b11111111111110100111, 
20'b11111111111101101000, 
20'b00000000000001111000, 
20'b11111111111110101000, 
20'b11111111111111001110, 
20'b11111111111101000001, 
20'b00000000000000100111, 
20'b11111111111110111001, 
20'b00000000000000111101, 
20'b11111111111110010110, 
20'b00000000000010100011, 
20'b11111111111101110011, 
20'b00000000000010100011, 
20'b11111111111110110101, 
20'b11111111111010011010, 
20'b00000000000000110011, 
20'b00000000000010011010, 
20'b00000000000000001011, 
20'b00000000000000011011, 
20'b00000000000000100001, 
20'b00000000000010100101, 
20'b11111111111110011100, 
20'b00000000000000101111, 
20'b11111111111100000111, 
20'b00000000000010000001, 
20'b00000000000010010001, 
20'b00000000000000010011, 
20'b11111111111110111100, 
20'b00000000000001010011, 
20'b11111111111111000010, 
20'b00000000000001000101, 
20'b00000000000000100011, 
20'b00000000000000000001, 
20'b00000000000000011000, 
20'b11111111111101100111, 
20'b00000000000000110000, 
20'b11111111111111010011, 
20'b00000000000000100111, 
20'b00000000000011010100, 
20'b00000000000010001011, 
20'b11111111111111101001, 
20'b11111111111100110101, 
20'b00000000000001110010, 
20'b11111111111100010101, 
20'b11111111111110111111, 
20'b11111111111110011110, 
20'b11111111111111111011, 
20'b00000000000010101111, 
20'b11111111111111001011, 
20'b00000000000000000010, 
20'b00000000000011111000, 
20'b11111111111111010001, 
20'b11111111111111010001, 
20'b11111111111110111100, 
20'b11111111111111101100, 
20'b00000000000010000100, 
20'b11111111111101001000, 
20'b11111111111110100111, 
20'b11111111111110101010, 
20'b11111111111100111010, 
20'b11111111111101111000, 
20'b11111111111011110100, 
20'b11111111111110010110, 
20'b11111111111110011100, 
20'b11111111111011111111, 
20'b00000000000011000110, 
20'b11111111111100111111, 
20'b00000000000001000110, 
20'b11111111111101010111, 
20'b11111111111101011001, 
20'b00000000000001111011, 
20'b00000000000000000011, 
20'b11111111111101001010, 
20'b00000000000000101110, 
20'b11111111111100101110, 
20'b00000000000010100100, 
20'b00000000000001001000, 
20'b11111111111110110100, 
20'b11111111111101111011, 
20'b11111111111110000011, 
20'b00000000000001100111, 
20'b11111111111101000000, 
20'b00000000000000001010, 
20'b00000000000010100100, 
20'b00000000000001011000, 
20'b00000000000001101101, 
20'b11111111111101001100, 
20'b00000000000011001111, 
20'b00000000000010011101, 
20'b00000000000000011001, 
20'b00000000000011101000, 
20'b00000000000000011101, 
20'b11111111111011100111, 
20'b00000000000011011000, 
20'b00000000000001010011, 
20'b00000000000010110011, 
20'b11111111111100011100, 
20'b11111111111111010011, 
20'b00000000000000111001, 
20'b11111111111101001110, 
20'b11111111111101100100, 
20'b11111111111101101110, 
20'b11111111111110010111, 
20'b00000000000011101010, 
20'b00000000000000001101, 
20'b00000000000001101000, 
20'b00000000000000001100, 
20'b00000000000011000010, 
20'b00000000000010111000, 
20'b11111111111100001111, 
20'b11111111111101011000, 
20'b00000000000010001101, 
20'b11111111111101111011, 
20'b11111111111111011000, 
20'b11111111111111011000, 
20'b00000000000010000011, 
20'b00000000000000110001, 
20'b11111111111111110111, 
20'b11111111111101010101, 
20'b00000000000010011110, 
20'b11111111111111001010, 
20'b00000000000010101110, 
20'b00000000000000111101, 
20'b00000000000001010101, 
20'b11111111111110111110, 
20'b00000000000000010001, 
20'b00000000000010101110, 
20'b11111111111111011101, 
20'b11111111111111110100, 
20'b11111111111111101000, 
20'b11111111111101100111, 
20'b00000000000100000001, 
20'b00000000000000100110, 
20'b11111111111110000101, 
20'b11111111111111101010, 
20'b00000000000000111000, 
20'b11111111111111010011, 
20'b11111111111111010001, 
20'b00000000000000100100, 
20'b00000000000011001011, 
20'b00000000000001110001, 
20'b00000000000010110110, 
20'b00000000000000111111, 
20'b11111111111101101000, 
20'b00000000000000101000, 
20'b11111111111101101000, 
20'b11111111111110101010, 
20'b11111111111110000100, 
20'b00000000000000000001, 
20'b00000000000000010110, 
20'b00000000000001010111, 
20'b00000000000000110011, 
20'b00000000000001000001, 
20'b11111111111011001110, 
20'b11111111111101100000, 
20'b11111111111111100001, 
20'b00000000000000011100, 
20'b00000000000011110110, 
20'b00000000000011110001, 
20'b11111111111011110011, 
20'b11111111111111011111, 
20'b00000000000010000100, 
20'b00000000000011010110, 
20'b11111111111011110011, 
20'b11111111111101101001, 
20'b00000000000000011100, 
20'b00000000000010010110, 
20'b11111111111110100011, 
20'b11111111111110111011, 
20'b11111111111111001001, 
20'b11111111111111110101, 
20'b00000000000011010110, 
20'b00000000000010101001, 
20'b11111111111111101101, 
20'b11111111111110110110, 
20'b00000000000010010110, 
20'b00000000000001001000, 
20'b00000000000010001010, 
20'b11111111111111100111, 
20'b11111111111110000111, 
20'b11111111111111000110, 
20'b11111111111111100100, 
20'b11111111111100101000, 
20'b00000000000000101101, 
20'b11111111111100110000, 
20'b00000000000001100111, 
20'b11111111111111100001, 
20'b11111111111111100101, 
20'b00000000000010000011, 
20'b00000000000000010011, 
20'b11111111111111101011, 
20'b00000000000001010110, 
20'b00000000000001000011, 
20'b00000000000000110111, 
20'b00000000000000011011, 
20'b00000000000001100000, 
20'b11111111111101111101, 
20'b00000000000100000010, 
20'b00000000000001111110, 
20'b11111111111011101001, 
20'b00000000000000010010, 
20'b11111111111100100001, 
20'b11111111111100011000, 
20'b11111111111011010111, 
20'b11111111111111001010, 
20'b11111111111110101011, 
20'b11111111111110000011, 
20'b00000000000001011011, 
20'b00000000000000010000, 
20'b11111111111100111110, 
20'b00000000000000101001, 
20'b11111111111110000110, 
20'b11111111111110010000, 
20'b11111111111110100000, 
20'b11111111111110111101, 
20'b11111111111110011000, 
20'b00000000000000010001, 
20'b11111111111111001001, 
20'b00000000000010010110, 
20'b11111111111110000001, 
20'b00000000000000110110, 
20'b00000000000000011001, 
20'b00000000000001011001, 
20'b00000000000011011001, 
20'b00000000000000000001, 
20'b11111111111101110101, 
20'b11111111111110100000, 
20'b00000000000001110010, 
20'b00000000000010001110, 
20'b11111111111010111101, 
20'b00000000000001001101, 
20'b00000000000000010011, 
20'b11111111111011101010, 
20'b00000000000010110101, 
20'b11111111111110110001, 
20'b00000000000000000100, 
20'b11111111111101101110, 
20'b00000000000010110000, 
20'b00000000000001111100, 
20'b11111111111010011010, 
20'b00000000000010001110, 
20'b00000000000001011111, 
20'b00000000000001011001, 
20'b00000000000100101001, 
20'b00000000000001010011, 
20'b00000000000010100010, 
20'b11111111111101100011, 
20'b00000000000000100100, 
20'b11111111111111000100, 
20'b00000000000001000100, 
20'b00000000000011101100, 
20'b00000000000001110110, 
20'b11111111111010111010, 
20'b00000000000010100110, 
20'b11111111111110110110, 
20'b00000000000000101101, 
20'b11111111111101111101, 
20'b11111111111101001001, 
20'b00000000000000100011, 
20'b00000000000001111000, 
20'b00000000000000111101, 
20'b11111111111111000110, 
20'b11111111111011011000, 
20'b00000000000001001010, 
20'b00000000000000011011, 
20'b00000000000010010100, 
20'b00000000000000000110, 
20'b00000000000000100010, 
20'b00000000000010011101, 
20'b00000000000010001000, 
20'b11111111111110110110, 
20'b00000000000001101110, 
20'b11111111111101111101, 
20'b11111111111101111110, 
20'b11111111111110101000, 
20'b00000000000010110010, 
20'b11111111111110000111, 
20'b11111111111101001111, 
20'b00000000000000011101, 
20'b00000000000001101111, 
20'b00000000000010001001, 
20'b11111111111110011101, 
20'b11111111111011101110, 
20'b11111111111011100111, 
20'b00000000000001111010, 
20'b00000000000000001111, 
20'b00000000000010101110, 
20'b00000000000010001101, 
20'b00000000000001110111, 
20'b00000000000010111000, 
20'b11111111111110100111, 
20'b11111111111111110000, 
20'b00000000000000101101, 
20'b00000000000001001010, 
20'b00000000000010011100, 
20'b00000000000010101110, 
20'b00000000000011010000, 
20'b11111111111101111001, 
20'b00000000000000000001, 
20'b00000000000011010100, 
20'b00000000000010011011, 
20'b00000000000010010001, 
20'b11111111111111110011, 
20'b11111111111101011111, 
20'b11111111111111010100, 
20'b11111111111111011010, 
20'b11111111111101111000, 
20'b11111111111100000100, 
20'b00000000000010000111, 
20'b00000000000001111000, 
20'b00000000000010100001, 
20'b00000000000000000010, 
20'b11111111111110011110, 
20'b11111111111111010111, 
20'b11111111111110000110, 
20'b00000000000000011110, 
20'b00000000000000000010, 
20'b00000000000010111101, 
20'b00000000000001010011, 
20'b11111111111011100010, 
20'b11111111111101101110, 
20'b11111111111101001011, 
20'b11111111111111111001, 
20'b11111111111100011000, 
20'b11111111111111001111, 
20'b11111111111110110100, 
20'b00000000000000110111, 
20'b00000000000000001001, 
20'b00000000000000100011, 
20'b11111111111011001101, 
20'b11111111111111110100, 
20'b00000000000010001010, 
20'b00000000000011011000, 
20'b11111111111111101010, 
20'b11111111111100001111, 
20'b00000000000001111001, 
20'b11111111111111000110, 
20'b00000000000010110101, 
20'b11111111111111111010, 
20'b11111111111011011111, 
20'b11111111111110100001, 
20'b00000000000000010110, 
20'b11111111111100010011, 
20'b11111111111111101010, 
20'b00000000000010110100, 
20'b11111111111110110100, 
20'b11111111111111110101, 
20'b00000000000010101111, 
20'b00000000000000111011, 
20'b11111111111110110111, 
20'b00000000000010111000, 
20'b11111111111110111000, 
20'b00000000000001001100, 
20'b00000000000000001101, 
20'b11111111111100111010, 
20'b00000000000010100001, 
20'b11111111111110011011, 
20'b00000000000000001001, 
20'b00000000000000010100, 
20'b11111111111110100111, 
20'b11111111111111001100, 
20'b00000000000001110001, 
20'b00000000000000000010, 
20'b00000000000000101101, 
20'b00000000000001001101, 
20'b11111111111110001110, 
20'b00000000000000111010, 
20'b11111111111101010110, 
20'b11111111111111111011, 
20'b11111111111110011011, 
20'b11111111111110010100, 
20'b11111111111101100100, 
20'b00000000000000011000, 
20'b00000000000001010100, 
20'b00000000000000101111, 
20'b11111111111110110000, 
20'b11111111111101101010, 
20'b00000000000010101001, 
20'b11111111111110011111, 
20'b00000000000000000001, 
20'b00000000000011001111, 
20'b00000000000000000100, 
20'b11111111111100110010, 
20'b00000000000010001101, 
20'b11111111111101110011, 
20'b00000000000001011101, 
20'b00000000000000111111, 
20'b00000000000001000001, 
20'b00000000000010000111, 
20'b11111111111101100001, 
20'b00000000000000110010, 
20'b11111111111110011000, 
20'b11111111111101000101, 
20'b00000000000001101110, 
20'b11111111111100111010, 
20'b00000000000010110101, 
20'b00000000000000100010, 
20'b11111111111110111000, 
20'b11111111111100110010, 
20'b11111111111110100111, 
20'b00000000000010101001, 
20'b11111111111110000011, 
20'b00000000000000001010, 
20'b11111111111110101001, 
20'b00000000000011000000, 
20'b11111111111111011110, 
20'b00000000000000010011, 
20'b00000000000001100001, 
20'b11111111111110011010, 
20'b11111111111110001100, 
20'b00000000000000110000, 
20'b00000000000000011001, 
20'b11111111111100010100, 
20'b00000000000011011010, 
20'b11111111111111010010, 
20'b00000000000011001010, 
20'b00000000000001110001, 
20'b00000000000001100100, 
20'b11111111111101110000, 
20'b11111111111111010000, 
20'b11111111111111010000, 
20'b11111111111110111000, 
20'b11111111111111101011, 
20'b00000000000001110001, 
20'b11111111111110000011, 
20'b00000000000001100110, 
20'b00000000000000010111, 
20'b00000000000000100010, 
20'b00000000000001101001, 
20'b00000000000010100001, 
20'b00000000000001010101, 
20'b11111111111110001000, 
20'b00000000000000111010, 
20'b11111111111100001111, 
20'b00000000000001000100, 
20'b11111111111110110100, 
20'b00000000000001100010, 
20'b11111111111110100100, 
20'b11111111111110010011, 
20'b00000000000001010101, 
20'b11111111111101100011, 
20'b11111111111110011111, 
20'b11111111111101010011, 
20'b00000000000000011101, 
20'b11111111111110001101, 
20'b00000000000011100110, 
20'b11111111111111101001, 
20'b11111111111110001000, 
20'b11111111111111111100, 
20'b00000000000001010010, 
20'b00000000000001010000, 
20'b00000000000010101111, 
20'b11111111111110101111, 
20'b11111111111101000000, 
20'b00000000000000001101, 
20'b11111111111101111011, 
20'b11111111111110101110, 
20'b11111111111100100000, 
20'b00000000000001101100, 
20'b00000000000100001101, 
20'b00000000000001100111, 
20'b00000000000010100111, 
20'b11111111111111111001, 
20'b11111111111110001100, 
20'b00000000000010010000, 
20'b11111111111111000011, 
20'b00000000000010100011, 
20'b11111111111110110011, 
20'b00000000000000101110, 
20'b11111111111101000110, 
20'b00000000000100011000, 
20'b00000000000011110010, 
20'b11111111111110010011, 
20'b11111111111010111001, 
20'b00000000000000010111, 
20'b11111111111101100011, 
20'b00000000000100000011, 
20'b11111111111111100000, 
20'b11111111111110011011, 
20'b00000000000000011010, 
20'b11111111111110001100, 
20'b11111111111110010101, 
20'b11111111111110111011, 
20'b11111111111011001111, 
20'b00000000000000011110, 
20'b11111111111011010100, 
20'b11111111111110101010, 
20'b00000000000000011011, 
20'b00000000000001011101, 
20'b11111111111110001111, 
20'b11111111111111101110, 
20'b00000000000000101000, 
20'b11111111111110110110, 
20'b11111111111010101000, 
20'b11111111111110110101, 
20'b00000000000000110101, 
20'b00000000000000100101, 
20'b00000000000001001010, 
20'b00000000000001010001, 
20'b11111111111011101110, 
20'b11111111111110100000, 
20'b00000000000010110001, 
20'b11111111111100111001, 
20'b11111111111110111000, 
20'b00000000000011101110, 
20'b11111111111110011000, 
20'b00000000000000000110, 
20'b11111111111110011100, 
20'b00000000000000100001, 
20'b11111111111111010111, 
20'b11111111111110111001, 
20'b00000000000010111110, 
20'b11111111111100111111, 
20'b11111111111110111001, 
20'b00000000000010010010, 
20'b00000000000010111010, 
20'b11111111111111001010, 
20'b00000000000001000010, 
20'b11111111111111011000, 
20'b11111111111011101000, 
20'b11111111111110111100, 
20'b00000000000000100100, 
20'b11111111111110011100, 
20'b11111111111111111000, 
20'b11111111111111000000, 
20'b11111111111110011100, 
20'b00000000000010011010, 
20'b11111111111110011101, 
20'b11111111111110000000, 
20'b00000000000000001100, 
20'b11111111111111000000, 
20'b00000000000001010001, 
20'b11111111111101011000, 
20'b00000000000010100000, 
20'b00000000000001111111, 
20'b00000000000000001011, 
20'b11111111111111111010, 
20'b11111111111101110001, 
20'b11111111111101010110, 
20'b11111111111110001100, 
20'b11111111111110110110, 
20'b11111111111111011110, 
20'b00000000000000101000, 
20'b00000000000011110011, 
20'b11111111111110111010, 
20'b11111111111100011101, 
20'b00000000000011101011, 
20'b11111111111110001101, 
20'b11111111111111100100, 
20'b00000000000000100010, 
20'b00000000000001101011, 
20'b11111111111101111101, 
20'b11111111111110001000, 
20'b11111111111111001100, 
20'b00000000000001110111, 
20'b11111111111110011101, 
20'b00000000000001100101, 
20'b00000000000001110101, 
20'b11111111111101001100, 
20'b00000000000000000111, 
20'b00000000000000000011, 
20'b11111111111111001100, 
20'b11111111111110110010, 
20'b00000000000000010110, 
20'b11111111111111001110, 
20'b00000000000000111001, 
20'b00000000000000110110, 
20'b11111111111101010010, 
20'b11111111111110001001, 
20'b00000000000000011101, 
20'b00000000000001111000, 
20'b11111111111100100001, 
20'b11111111111011100111, 
20'b11111111111110011100, 
20'b11111111111111010011, 
20'b11111111111111011110, 
20'b11111111111111101101, 
20'b11111111111101101101, 
20'b00000000000001010110, 
20'b00000000000001011110, 
20'b11111111111110011101, 
20'b00000000000001101101, 
20'b11111111111111110001, 
20'b11111111111110111010, 
20'b00000000000010110001, 
20'b11111111111110000111, 
20'b11111111111111011011, 
20'b11111111111110000110, 
20'b00000000000000110010, 
20'b00000000000010010001, 
20'b11111111111111111000, 
20'b00000000000001011011, 
20'b11111111111011011100, 
20'b00000000000000011011, 
20'b11111111111110010111, 
20'b11111111111110101100, 
20'b00000000000010011010, 
20'b11111111111101000111, 
20'b00000000000001010100, 
20'b11111111111110101111, 
20'b00000000000000000100, 
20'b00000000000000000100, 
20'b11111111111100110010, 
20'b11111111111111110011, 
20'b00000000000000011110, 
20'b11111111111101101101, 
20'b00000000000000100000, 
20'b00000000000010100000, 
20'b11111111111110010001, 
20'b00000000000001111001, 
20'b11111111111111000111, 
20'b00000000000011011110, 
20'b11111111111010111110, 
20'b11111111111010110001, 
20'b00000000000001100011, 
20'b11111111111110100100, 
20'b00000000000000101010, 
20'b11111111111101110111, 
20'b11111111111111010111, 
20'b00000000000001110110, 
20'b00000000000000100010, 
20'b11111111111111111000, 
20'b00000000000000100000, 
20'b11111111111110010010, 
20'b00000000000010001011, 
20'b11111111111111111011, 
20'b11111111111110011101, 
20'b00000000000001010001, 
20'b11111111111111100010, 
20'b00000000000000001110, 
20'b00000000000001111101, 
20'b11111111111100100111, 
20'b11111111111110000001, 
20'b11111111111010111101, 
20'b00000000000001000000, 
20'b11111111111100100101, 
20'b00000000000001100000, 
20'b00000000000001001111, 
20'b11111111111111111111, 
20'b11111111111101111110, 
20'b11111111111110010111, 
20'b00000000000001110011, 
20'b11111111111111101001, 
20'b11111111111011111100, 
20'b00000000000011001011, 
20'b11111111111011100010, 
20'b11111111111101100110, 
20'b11111111111111100001, 
20'b00000000000000000001, 
20'b11111111111101001001, 
20'b11111111111110101101, 
20'b11111111111111111100, 
20'b11111111111111101101, 
20'b11111111111111010000, 
20'b11111111111111110101, 
20'b11111111111110001011, 
20'b00000000000011100011, 
20'b11111111111111000100, 
20'b00000000000000011100, 
20'b00000000000000011101, 
20'b11111111111111011000, 
20'b00000000000000101001, 
20'b00000000000000010111, 
20'b11111111111111001111, 
20'b11111111111111010011, 
20'b00000000000000110110, 
20'b00000000000000011010, 
20'b00000000000000101100, 
20'b00000000000001010110, 
20'b11111111111101101000, 
20'b00000000000011111001, 
20'b11111111111110100001, 
20'b00000000000000100001, 
20'b11111111111110101000, 
20'b00000000000001010011, 
20'b11111111111101001110, 
20'b11111111111101110011, 
20'b11111111111100011101, 
20'b11111111111111010100, 
20'b11111111111010110010, 
20'b11111111111111110110, 
20'b11111111111110001111, 
20'b11111111111101001000, 
20'b11111111111101111000, 
20'b11111111111110111110, 
20'b11111111111110001000, 
20'b00000000000010101000, 
20'b11111111111010111101, 
20'b00000000000100001000, 
20'b11111111111111010111, 
20'b11111111111101111011, 
20'b11111111111111010101, 
20'b11111111111100111011, 
20'b00000000000000100100, 
20'b00000000000001011000, 
20'b11111111111101010110, 
20'b00000000000000101110, 
20'b11111111111100010010, 
20'b00000000000010000100, 
20'b11111111111100111111, 
20'b00000000000000101111, 
20'b11111111111110100010, 
20'b11111111111111000011, 
20'b00000000000010110010, 
20'b00000000000010010010, 
20'b11111111111110011000, 
20'b00000000000010001111, 
20'b00000000000000111000, 
20'b00000000000000100110, 
20'b00000000000011011010, 
20'b00000000000001111101, 
20'b11111111111110010000, 
20'b11111111111110000001, 
20'b00000000000010111000, 
20'b00000000000010101011, 
20'b00000000000000001110, 
20'b00000000000001100001, 
20'b00000000000000101111, 
20'b00000000000000101101, 
20'b11111111111111011000, 
20'b00000000000010011110, 
20'b11111111111111100001, 
20'b00000000000000000011, 
20'b00000000000000111101, 
20'b00000000000100110010, 
20'b11111111111101010110, 
20'b11111111111110111011, 
20'b00000000000000000111, 
20'b00000000000010000000, 
20'b00000000000010011111, 
20'b11111111111101100011, 
20'b11111111111101011000, 
20'b00000000000000010100, 
20'b00000000000000111001, 
20'b00000000000000010100, 
20'b00000000000000100001, 
20'b00000000000001001000, 
20'b00000000000000111010, 
20'b00000000000010000100, 
20'b11111111111111111001, 
20'b00000000000000010110, 
20'b00000000000010010000, 
20'b11111111111111110110, 
20'b11111111111111010001, 
20'b00000000000000100001, 
20'b11111111111100110011, 
20'b00000000000000011000, 
20'b00000000000001011001, 
20'b11111111111101011101, 
20'b00000000000011111011, 
20'b11111111111111110001, 
20'b00000000000000111110, 
20'b11111111111111110101, 
20'b11111111111111011011, 
20'b11111111111111010010, 
20'b00000000000001110111, 
20'b00000000000011111100, 
20'b00000000000000000000, 
20'b00000000000001100001, 
20'b00000000000100000010, 
20'b11111111111100111100, 
20'b00000000000001111000, 
20'b00000000000010000011, 
20'b11111111111101111011, 
20'b00000000000000011111, 
20'b00000000000010011101, 
20'b00000000000000001111, 
20'b00000000000001110100, 
20'b11111111111111101110, 
20'b00000000000011011100, 
20'b00000000000001011110, 
20'b11111111111110100011, 
20'b11111111111100001110, 
20'b11111111111101101110, 
20'b00000000000000110010, 
20'b00000000000000001110, 
20'b11111111111111100001, 
20'b00000000000001000111, 
20'b00000000000001011010, 
20'b00000000000001010100, 
20'b11111111111100011001, 
20'b00000000000000101111, 
20'b00000000000001101001, 
20'b11111111111100110110, 
20'b11111111111110010111, 
20'b11111111111111011101, 
20'b00000000000011001001, 
20'b00000000000011010101, 
20'b11111111111111111100, 
20'b00000000000001110101, 
20'b11111111111100110101, 
20'b11111111111110110101, 
20'b11111111111110111100, 
20'b11111111111111100101, 
20'b00000000000000010010, 
20'b11111111111011110000, 
20'b00000000000001110110, 
20'b11111111111111001011, 
20'b11111111111111001000, 
20'b11111111111101010000, 
20'b00000000000000011101, 
20'b11111111111111110111, 
20'b00000000000100101111, 
20'b11111111111100010111, 
20'b00000000000001000000, 
20'b00000000000000000111, 
20'b11111111111110000101, 
20'b11111111111110110010, 
20'b00000000000000101001, 
20'b11111111111101010110, 
20'b11111111111110011101, 
20'b11111111111100011110, 
20'b11111111111111000110, 
20'b00000000000001101110, 
20'b00000000000011001100, 
20'b11111111111101111011, 
20'b11111111111111001100, 
20'b00000000000000100110, 
20'b00000000000010100101, 
20'b11111111111110111101, 
20'b11111111111111111100, 
20'b11111111111111101010, 
20'b00000000000010110001, 
20'b11111111111011101110, 
20'b00000000000010101011, 
20'b11111111111110010000, 
20'b11111111111011111001, 
20'b11111111111101111000, 
20'b00000000000100001010, 
20'b11111111111100101110, 
20'b11111111111111000100, 
20'b11111111111100000010, 
20'b00000000000001100011, 
20'b00000000000011100001, 
20'b00000000000011101100, 
20'b11111111111101111100, 
20'b00000000000000001100, 
20'b11111111111011110010, 
20'b00000000000001101101, 
20'b11111111111110000100, 
20'b00000000000010010111, 
20'b00000000000000000101, 
20'b00000000000001010000, 
20'b11111111111110000010, 
20'b11111111111110011011, 
20'b11111111111101110111, 
20'b00000000000000110011, 
20'b00000000000001000110, 
20'b00000000000011011111, 
20'b00000000000000100010, 
20'b11111111111110000101, 
20'b11111111111111000011, 
20'b11111111111100100100, 
20'b00000000000010101010, 
20'b00000000000001110110, 
20'b11111111111101000100, 
20'b11111111111111001110, 
20'b11111111111011110011, 
20'b00000000000010101011, 
20'b11111111111100110010, 
20'b00000000000011010001, 
20'b11111111111101111110, 
20'b00000000000000110001, 
20'b00000000000000011011, 
20'b00000000000010100001, 
20'b11111111111101101111, 
20'b11111111111101011111, 
20'b00000000000010110100, 
20'b11111111111110011011, 
20'b00000000000000010100, 
20'b11111111111101010100, 
20'b00000000000000001100, 
20'b11111111111110100001, 
20'b00000000000001110101, 
20'b11111111111110110101, 
20'b11111111111110011010, 
20'b11111111111110100001, 
20'b00000000000001100100, 
20'b11111111111110110010, 
20'b11111111111111010101, 
20'b00000000000001010001, 
20'b00000000000010011011, 
20'b11111111111100001011, 
20'b00000000000000010010, 
20'b00000000000000011011, 
20'b11111111111011111001, 
20'b11111111111111011001, 
20'b00000000000011000101, 
20'b00000000000001110100, 
20'b11111111111100011101, 
20'b00000000000001111011, 
20'b11111111111001000100, 
20'b11111111111100101111, 
20'b11111111111101001010, 
20'b00000000000000010000, 
20'b11111111111011101010, 
20'b11111111111110111001, 
20'b00000000000000010010, 
20'b11111111111110100000, 
20'b00000000000011111111, 
20'b00000000000000100000, 
20'b00000000000000001010, 
20'b00000000000000000000, 
20'b00000000000100101100, 
20'b11111111111101001110, 
20'b11111111111101011111, 
20'b00000000000000101110, 
20'b00000000000010101000, 
20'b00000000000010000001, 
20'b00000000000010000011, 
20'b11111111111110001010, 
20'b11111111111101011110, 
20'b00000000000000011110, 
20'b11111111111101110101, 
20'b00000000000000101011, 
20'b00000000000000111110, 
20'b00000000000000010100, 
20'b11111111111100010111, 
20'b11111111111100010101, 
20'b11111111111111100100, 
20'b11111111111111000111, 
20'b11111111111111011011, 
20'b11111111111100000101, 
20'b00000000000000101011, 
20'b11111111111110101001, 
20'b11111111111011010101, 
20'b11111111111101111010, 
20'b00000000000010101110, 
20'b11111111111100111101, 
20'b00000000000010010011, 
20'b00000000000100000010, 
20'b00000000000011111100, 
20'b11111111111111111000, 
20'b11111111111101010111, 
20'b00000000000001101111, 
20'b11111111111101011000, 
20'b11111111111110111000, 
20'b00000000000001100111, 
20'b11111111111111100100, 
20'b11111111111111011111, 
20'b11111111111111011011, 
20'b00000000000010000011

};
localparam logic signed [19:0] dlBiases [9:0] = {
20'b00000000000010101010, 
20'b11111111111111111110, 
20'b11111111111111111110, 
20'b11111111111111000100, 
20'b11111111111111000001, 
20'b11111111111111101011, 
20'b11111111111111101001, 
20'b00000000000001001110, 
20'b11111111111101000111, 
20'b11111111111111101011

};
localparam logic signed [19:0] convWeights [0:17] = {
20'b00000000000001110010, 
20'b00000000000111101100, 
20'b11111111111100001011, 
20'b00000000000001011111, 
20'b00000000000000001110, 
20'b00000000001000001101, 
20'b00000000000110011111, 
20'b00000000000011001100, 
20'b11111111111100010110, 
20'b00000000000101100100, 
20'b11111111111110100111, 
20'b00000000000011010111, 
20'b00000000000111111101, 
20'b00000000000010100011, 
20'b00000000000110001000, 
20'b11111111111111110100, 
20'b00000000000010111010, 
20'b00000000000001110100 

};
localparam logic signed [19:0] convBiases [1:0] = {
20'b00000000000000000000, 
20'b00000000000000000000

};
endpackage