package data4_2;

localparam logic signed [3:0] dlWeights [0:1279] = {
4'b0001, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0001, 
4'b0010, 
4'b1110, 
4'b1111, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0001, 
4'b1111, 
4'b1110, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b1111, 
4'b0001, 
4'b1110, 
4'b1110, 
4'b0000, 
4'b0001, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1110, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0001, 
4'b1111, 
4'b1110, 
4'b1111, 
4'b0001, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1110, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1100, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1110, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0001, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1110, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1110, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0001, 
4'b1110, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1110, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b0000, 
4'b0000, 
4'b0001, 
4'b1110, 
4'b1111, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1110, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1110, 
4'b1111, 
4'b1111, 
4'b1110, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0001, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0001, 
4'b0000, 
4'b1110, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1110, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0001, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1110, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1110, 
4'b1110, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0001, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0001, 
4'b0000, 
4'b1111, 
4'b1110, 
4'b0000, 
4'b1111, 
4'b0001, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1110, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1110, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1110, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1110, 
4'b1110, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1110, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1110, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1110, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1110, 
4'b0001, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0001, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0001, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1110, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0001, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1110, 
4'b0000, 
4'b1111, 
4'b1110, 
4'b1111, 
4'b0001, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1110, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1110, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0001, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1110, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b0000, 
4'b0001, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000
};
localparam logic signed [3:0] dlBiases [9:0] = {
4'b0000, 
4'b0000, 
4'b0000, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b1111, 
4'b0000, 
4'b1111, 
4'b1111
};
localparam logic signed [3:0] convWeights [0:17] = {
4'b0000, 
4'b0001, 
4'b1111, 
4'b0000, 
4'b0000, 
4'b0010, 
4'b0001, 
4'b0000, 
4'b1111, 
4'b0001, 
4'b1111, 
4'b0000, 
4'b0001, 
4'b0000, 
4'b0001, 
4'b1111, 
4'b0000, 
4'b0000
};

localparam logic signed [3:0] convBiases [1:0] = {
4'b0000, 
4'b0000 
};

endpackage