package data8_4;
localparam logic signed [7:0] dlWeights [0:1279] = {
8'b00000100, 
8'b00000000, 
8'b11111100, 
8'b00000000, 
8'b11111110, 
8'b00000010, 
8'b00000001, 
8'b11111100, 
8'b00000000, 
8'b00000010, 
8'b00000010, 
8'b11111011, 
8'b11111001, 
8'b11111101, 
8'b00000001, 
8'b11111110, 
8'b11111110, 
8'b11111111, 
8'b11111111, 
8'b11111111, 
8'b00000001, 
8'b11111100, 
8'b00000000, 
8'b00000001, 
8'b11111111, 
8'b00000000, 
8'b11111110, 
8'b00000000, 
8'b00000001, 
8'b00000100, 
8'b00001001, 
8'b11111001, 
8'b11111100, 
8'b11111011, 
8'b11111100, 
8'b00000001, 
8'b11111111, 
8'b00000010, 
8'b11111110, 
8'b00000011, 
8'b00000010, 
8'b11111101, 
8'b11111111, 
8'b11111101, 
8'b00000000, 
8'b11111110, 
8'b00000010, 
8'b11111101, 
8'b11111110, 
8'b00000000, 
8'b00000101, 
8'b11111101, 
8'b11111011, 
8'b11111010, 
8'b11111101, 
8'b00000001, 
8'b11111111, 
8'b00000010, 
8'b00000001, 
8'b00000001, 
8'b00000011, 
8'b11111100, 
8'b00000001, 
8'b00000001, 
8'b11111101, 
8'b00000011, 
8'b00000011, 
8'b00000000, 
8'b00000010, 
8'b11111110, 
8'b00000000, 
8'b00000011, 
8'b11111100, 
8'b11111101, 
8'b11111101, 
8'b00000001, 
8'b11111111, 
8'b00000010, 
8'b11111100, 
8'b11111101, 
8'b11111110, 
8'b11111110, 
8'b11111100, 
8'b00000001, 
8'b11111101, 
8'b00000010, 
8'b00000000, 
8'b11111101, 
8'b11111111, 
8'b11111110, 
8'b00000000, 
8'b00000000, 
8'b11111110, 
8'b00000000, 
8'b11111011, 
8'b11111111, 
8'b11111100, 
8'b00000101, 
8'b11111011, 
8'b11111011, 
8'b00000000, 
8'b00000100, 
8'b00000000, 
8'b00000000, 
8'b11111101, 
8'b11111111, 
8'b11111101, 
8'b11111101, 
8'b00000001, 
8'b11111100, 
8'b00000000, 
8'b00000010, 
8'b00000000, 
8'b00000010, 
8'b11111100, 
8'b11111110, 
8'b11111011, 
8'b00000001, 
8'b11111101, 
8'b00000001, 
8'b11111101, 
8'b11111111, 
8'b00000000, 
8'b00000001, 
8'b11111100, 
8'b11111110, 
8'b11111100, 
8'b11111110, 
8'b00000000, 
8'b00000001, 
8'b11111101, 
8'b11111110, 
8'b11111110, 
8'b00000100, 
8'b11111101, 
8'b11111010, 
8'b11111101, 
8'b00000101, 
8'b11111111, 
8'b00000000, 
8'b11111111, 
8'b11111110, 
8'b00000000, 
8'b00000000, 
8'b00000011, 
8'b11111111, 
8'b11111011, 
8'b00000011, 
8'b11111111, 
8'b00000001, 
8'b00000000, 
8'b00000001, 
8'b00000010, 
8'b11111111, 
8'b00000001, 
8'b11111101, 
8'b11110011, 
8'b00000011, 
8'b11111111, 
8'b00000001, 
8'b00000010, 
8'b11111111, 
8'b11111011, 
8'b00000010, 
8'b00000011, 
8'b11111110, 
8'b00000100, 
8'b11111111, 
8'b00000000, 
8'b11111111, 
8'b00000010, 
8'b11111111, 
8'b11111111, 
8'b11111010, 
8'b00000000, 
8'b00000000, 
8'b11111110, 
8'b11111111, 
8'b11111110, 
8'b00000010, 
8'b00000011, 
8'b11111100, 
8'b11111111, 
8'b11111110, 
8'b00000011, 
8'b11111111, 
8'b00000010, 
8'b11111110, 
8'b00000011, 
8'b00000000, 
8'b00000011, 
8'b11111010, 
8'b11111101, 
8'b11111011, 
8'b11111111, 
8'b00000001, 
8'b00000000, 
8'b00000001, 
8'b00000010, 
8'b11111111, 
8'b00000011, 
8'b11111011, 
8'b11111110, 
8'b11111101, 
8'b11111111, 
8'b00000000, 
8'b00000000, 
8'b11111111, 
8'b00000000, 
8'b11111110, 
8'b11111111, 
8'b11111111, 
8'b11111111, 
8'b11111100, 
8'b11111111, 
8'b00000000, 
8'b00000011, 
8'b11111110, 
8'b00000000, 
8'b00000000, 
8'b11111101, 
8'b11111111, 
8'b11111100, 
8'b00000010, 
8'b11111100, 
8'b00000011, 
8'b11111101, 
8'b00000000, 
8'b11111110, 
8'b11111011, 
8'b00000010, 
8'b00000011, 
8'b11111100, 
8'b00000001, 
8'b11111111, 
8'b00000000, 
8'b11111110, 
8'b00000010, 
8'b00000000, 
8'b00000000, 
8'b00000000, 
8'b11111110, 
8'b00000001, 
8'b00000001, 
8'b00000001, 
8'b11111110, 
8'b11111101, 
8'b11111110, 
8'b00000001, 
8'b11111101, 
8'b00000001, 
8'b00000001, 
8'b11111110, 
8'b11111101, 
8'b11111011, 
8'b11111110, 
8'b00000000, 
8'b00000000, 
8'b11111011, 
8'b11111100, 
8'b11111100, 
8'b00000000, 
8'b00000000, 
8'b00000001, 
8'b11111010, 
8'b00000000, 
8'b00000001, 
8'b11111100, 
8'b00000000, 
8'b11111111, 
8'b00000000, 
8'b00000010, 
8'b00000000, 
8'b00000000, 
8'b11111111, 
8'b11111100, 
8'b11111100, 
8'b00000100, 
8'b11111011, 
8'b00000000, 
8'b11111111, 
8'b00000000, 
8'b00000001, 
8'b11111111, 
8'b00000000, 
8'b11111110, 
8'b00000001, 
8'b11111111, 
8'b00000010, 
8'b00000001, 
8'b11111110, 
8'b00000001, 
8'b00000001, 
8'b00000000, 
8'b00000001, 
8'b11111110, 
8'b11111011, 
8'b11111111, 
8'b11111101, 
8'b11111110, 
8'b00000000, 
8'b00000011, 
8'b00000000, 
8'b00000001, 
8'b11111110, 
8'b00000000, 
8'b00000001, 
8'b11111110, 
8'b00000001, 
8'b00000011, 
8'b00000001, 
8'b00000001, 
8'b11111111, 
8'b00000000, 
8'b00000010, 
8'b00000001, 
8'b11111100, 
8'b00000000, 
8'b11111111, 
8'b11111111, 
8'b00000010, 
8'b11111011, 
8'b11111101, 
8'b00000001, 
8'b00000011, 
8'b00000000, 
8'b00000011, 
8'b11111011, 
8'b00000000, 
8'b00000001, 
8'b00000100, 
8'b11111011, 
8'b11111110, 
8'b11111010, 
8'b11111111, 
8'b00000001, 
8'b11111101, 
8'b00000000, 
8'b11111110, 
8'b11111101, 
8'b00000001, 
8'b11111110, 
8'b11111111, 
8'b11111101, 
8'b00000000, 
8'b11111110, 
8'b00000000, 
8'b11111110, 
8'b00000010, 
8'b11111101, 
8'b00000010, 
8'b11111110, 
8'b11111010, 
8'b00000000, 
8'b00000010, 
8'b00000000, 
8'b00000000, 
8'b00000000, 
8'b00000010, 
8'b11111110, 
8'b00000000, 
8'b11111100, 
8'b00000010, 
8'b00000010, 
8'b00000000, 
8'b11111110, 
8'b00000001, 
8'b11111111, 
8'b00000001, 
8'b00000000, 
8'b00000000, 
8'b00000000, 
8'b11111101, 
8'b00000000, 
8'b11111111, 
8'b00000000, 
8'b00000011, 
8'b00000010, 
8'b11111111, 
8'b11111100, 
8'b00000001, 
8'b11111100, 
8'b11111110, 
8'b11111110, 
8'b11111111, 
8'b00000010, 
8'b11111111, 
8'b00000000, 
8'b00000011, 
8'b11111111, 
8'b11111111, 
8'b11111110, 
8'b11111111, 
8'b00000010, 
8'b11111101, 
8'b11111110, 
8'b11111110, 
8'b11111100, 
8'b11111101, 
8'b11111011, 
8'b11111110, 
8'b11111110, 
8'b11111011, 
8'b00000011, 
8'b11111100, 
8'b00000001, 
8'b11111101, 
8'b11111101, 
8'b00000001, 
8'b00000000, 
8'b11111101, 
8'b00000000, 
8'b11111100, 
8'b00000010, 
8'b00000001, 
8'b11111110, 
8'b11111101, 
8'b11111110, 
8'b00000001, 
8'b11111101, 
8'b00000000, 
8'b00000010, 
8'b00000001, 
8'b00000001, 
8'b11111101, 
8'b00000011, 
8'b00000010, 
8'b00000000, 
8'b00000011, 
8'b00000000, 
8'b11111011, 
8'b00000011, 
8'b00000001, 
8'b00000010, 
8'b11111100, 
8'b11111111, 
8'b00000000, 
8'b11111101, 
8'b11111101, 
8'b11111101, 
8'b11111110, 
8'b00000011, 
8'b00000000, 
8'b00000001, 
8'b00000000, 
8'b00000011, 
8'b00000010, 
8'b11111100, 
8'b11111101, 
8'b00000010, 
8'b11111101, 
8'b11111111, 
8'b11111111, 
8'b00000010, 
8'b00000000, 
8'b11111111, 
8'b11111101, 
8'b00000010, 
8'b11111111, 
8'b00000010, 
8'b00000000, 
8'b00000001, 
8'b11111110, 
8'b00000000, 
8'b00000010, 
8'b11111111, 
8'b11111111, 
8'b11111111, 
8'b11111101, 
8'b00000100, 
8'b00000000, 
8'b11111110, 
8'b11111111, 
8'b00000000, 
8'b11111111, 
8'b11111111, 
8'b00000000, 
8'b00000011, 
8'b00000001, 
8'b00000010, 
8'b00000000, 
8'b11111101, 
8'b00000000, 
8'b11111101, 
8'b11111110, 
8'b11111110, 
8'b00000000, 
8'b00000000, 
8'b00000001, 
8'b00000000, 
8'b00000001, 
8'b11111011, 
8'b11111101, 
8'b11111111, 
8'b00000000, 
8'b00000011, 
8'b00000011, 
8'b11111011, 
8'b11111111, 
8'b00000010, 
8'b00000011, 
8'b11111011, 
8'b11111101, 
8'b00000000, 
8'b00000010, 
8'b11111110, 
8'b11111110, 
8'b11111111, 
8'b11111111, 
8'b00000011, 
8'b00000010, 
8'b11111111, 
8'b11111110, 
8'b00000010, 
8'b00000001, 
8'b00000010, 
8'b11111111, 
8'b11111110, 
8'b11111111, 
8'b11111111, 
8'b11111100, 
8'b00000000, 
8'b11111100, 
8'b00000001, 
8'b11111111, 
8'b11111111, 
8'b00000010, 
8'b00000000, 
8'b11111111, 
8'b00000001, 
8'b00000001, 
8'b00000000, 
8'b00000000, 
8'b00000001, 
8'b11111101, 
8'b00000100, 
8'b00000001, 
8'b11111011, 
8'b00000000, 
8'b11111100, 
8'b11111100, 
8'b11111011, 
8'b11111111, 
8'b11111110, 
8'b11111110, 
8'b00000001, 
8'b00000000, 
8'b11111100, 
8'b00000000, 
8'b11111110, 
8'b11111110, 
8'b11111110, 
8'b11111110, 
8'b11111110, 
8'b00000000, 
8'b11111111, 
8'b00000010, 
8'b11111110, 
8'b00000000, 
8'b00000000, 
8'b00000001, 
8'b00000011, 
8'b00000000, 
8'b11111101, 
8'b11111110, 
8'b00000001, 
8'b00000010, 
8'b11111010, 
8'b00000001, 
8'b00000000, 
8'b11111011, 
8'b00000010, 
8'b11111110, 
8'b00000000, 
8'b11111101, 
8'b00000010, 
8'b00000001, 
8'b11111010, 
8'b00000010, 
8'b00000001, 
8'b00000001, 
8'b00000100, 
8'b00000001, 
8'b00000010, 
8'b11111101, 
8'b00000000, 
8'b11111111, 
8'b00000001, 
8'b00000011, 
8'b00000001, 
8'b11111010, 
8'b00000010, 
8'b11111110, 
8'b00000000, 
8'b11111101, 
8'b11111101, 
8'b00000000, 
8'b00000001, 
8'b00000000, 
8'b11111111, 
8'b11111011, 
8'b00000001, 
8'b00000000, 
8'b00000010, 
8'b00000000, 
8'b00000000, 
8'b00000010, 
8'b00000010, 
8'b11111110, 
8'b00000001, 
8'b11111101, 
8'b11111101, 
8'b11111110, 
8'b00000010, 
8'b11111110, 
8'b11111101, 
8'b00000000, 
8'b00000001, 
8'b00000010, 
8'b11111110, 
8'b11111011, 
8'b11111011, 
8'b00000001, 
8'b00000000, 
8'b00000010, 
8'b00000010, 
8'b00000001, 
8'b00000010, 
8'b11111110, 
8'b11111111, 
8'b00000000, 
8'b00000001, 
8'b00000010, 
8'b00000010, 
8'b00000011, 
8'b11111101, 
8'b00000000, 
8'b00000011, 
8'b00000010, 
8'b00000010, 
8'b11111111, 
8'b11111101, 
8'b11111111, 
8'b11111111, 
8'b11111101, 
8'b11111100, 
8'b00000010, 
8'b00000001, 
8'b00000010, 
8'b00000000, 
8'b11111110, 
8'b11111111, 
8'b11111110, 
8'b00000000, 
8'b00000000, 
8'b00000010, 
8'b00000001, 
8'b11111011, 
8'b11111101, 
8'b11111101, 
8'b11111111, 
8'b11111100, 
8'b11111111, 
8'b11111110, 
8'b00000000, 
8'b00000000, 
8'b00000000, 
8'b11111011, 
8'b11111111, 
8'b00000010, 
8'b00000011, 
8'b11111111, 
8'b11111100, 
8'b00000001, 
8'b11111111, 
8'b00000010, 
8'b11111111, 
8'b11111011, 
8'b11111110, 
8'b00000000, 
8'b11111100, 
8'b11111111, 
8'b00000010, 
8'b11111110, 
8'b11111111, 
8'b00000010, 
8'b00000000, 
8'b11111110, 
8'b00000010, 
8'b11111110, 
8'b00000001, 
8'b00000000, 
8'b11111100, 
8'b00000010, 
8'b11111110, 
8'b00000000, 
8'b00000000, 
8'b11111110, 
8'b11111111, 
8'b00000001, 
8'b00000000, 
8'b00000000, 
8'b00000001, 
8'b11111110, 
8'b00000000, 
8'b11111101, 
8'b11111111, 
8'b11111110, 
8'b11111110, 
8'b11111101, 
8'b00000000, 
8'b00000001, 
8'b00000000, 
8'b11111110, 
8'b11111101, 
8'b00000010, 
8'b11111110, 
8'b00000000, 
8'b00000011, 
8'b00000000, 
8'b11111100, 
8'b00000010, 
8'b11111101, 
8'b00000001, 
8'b00000000, 
8'b00000001, 
8'b00000010, 
8'b11111101, 
8'b00000000, 
8'b11111110, 
8'b11111101, 
8'b00000001, 
8'b11111100, 
8'b00000010, 
8'b00000000, 
8'b11111110, 
8'b11111100, 
8'b11111110, 
8'b00000010, 
8'b11111110, 
8'b00000000, 
8'b11111110, 
8'b00000011, 
8'b11111111, 
8'b00000000, 
8'b00000001, 
8'b11111110, 
8'b11111110, 
8'b00000000, 
8'b00000000, 
8'b11111100, 
8'b00000011, 
8'b11111111, 
8'b00000011, 
8'b00000001, 
8'b00000001, 
8'b11111101, 
8'b11111111, 
8'b11111111, 
8'b11111110, 
8'b11111111, 
8'b00000001, 
8'b11111110, 
8'b00000001, 
8'b00000000, 
8'b00000000, 
8'b00000001, 
8'b00000010, 
8'b00000001, 
8'b11111110, 
8'b00000000, 
8'b11111100, 
8'b00000001, 
8'b11111110, 
8'b00000001, 
8'b11111110, 
8'b11111110, 
8'b00000001, 
8'b11111101, 
8'b11111110, 
8'b11111101, 
8'b00000000, 
8'b11111110, 
8'b00000011, 
8'b11111111, 
8'b11111110, 
8'b11111111, 
8'b00000001, 
8'b00000001, 
8'b00000010, 
8'b11111110, 
8'b11111101, 
8'b00000000, 
8'b11111101, 
8'b11111110, 
8'b11111100, 
8'b00000001, 
8'b00000100, 
8'b00000001, 
8'b00000010, 
8'b11111111, 
8'b11111110, 
8'b00000010, 
8'b11111111, 
8'b00000010, 
8'b11111110, 
8'b00000000, 
8'b11111101, 
8'b00000100, 
8'b00000011, 
8'b11111110, 
8'b11111010, 
8'b00000000, 
8'b11111101, 
8'b00000100, 
8'b11111111, 
8'b11111110, 
8'b00000000, 
8'b11111110, 
8'b11111110, 
8'b11111110, 
8'b11111011, 
8'b00000000, 
8'b11111011, 
8'b11111110, 
8'b00000000, 
8'b00000001, 
8'b11111110, 
8'b11111111, 
8'b00000000, 
8'b11111110, 
8'b11111010, 
8'b11111110, 
8'b00000000, 
8'b00000000, 
8'b00000001, 
8'b00000001, 
8'b11111011, 
8'b11111110, 
8'b00000010, 
8'b11111100, 
8'b11111110, 
8'b00000011, 
8'b11111110, 
8'b00000000, 
8'b11111110, 
8'b00000000, 
8'b11111111, 
8'b11111110, 
8'b00000010, 
8'b11111100, 
8'b11111110, 
8'b00000010, 
8'b00000010, 
8'b11111111, 
8'b00000001, 
8'b11111111, 
8'b11111011, 
8'b11111110, 
8'b00000000, 
8'b11111110, 
8'b11111111, 
8'b11111111, 
8'b11111110, 
8'b00000010, 
8'b11111110, 
8'b11111110, 
8'b00000000, 
8'b11111111, 
8'b00000001, 
8'b11111101, 
8'b00000010, 
8'b00000001, 
8'b00000000, 
8'b11111111, 
8'b11111101, 
8'b11111101, 
8'b11111110, 
8'b11111110, 
8'b11111111, 
8'b00000000, 
8'b00000011, 
8'b11111110, 
8'b11111100, 
8'b00000011, 
8'b11111110, 
8'b11111111, 
8'b00000000, 
8'b00000001, 
8'b11111101, 
8'b11111110, 
8'b11111111, 
8'b00000001, 
8'b11111110, 
8'b00000001, 
8'b00000001, 
8'b11111101, 
8'b00000000, 
8'b00000000, 
8'b11111111, 
8'b11111110, 
8'b00000000, 
8'b11111111, 
8'b00000000, 
8'b00000000, 
8'b11111101, 
8'b11111110, 
8'b00000000, 
8'b00000001, 
8'b11111100, 
8'b11111011, 
8'b11111110, 
8'b11111111, 
8'b11111111, 
8'b11111111, 
8'b11111101, 
8'b00000001, 
8'b00000001, 
8'b11111110, 
8'b00000001, 
8'b11111111, 
8'b11111110, 
8'b00000010, 
8'b11111110, 
8'b11111111, 
8'b11111110, 
8'b00000000, 
8'b00000010, 
8'b11111111, 
8'b00000001, 
8'b11111011, 
8'b00000000, 
8'b11111110, 
8'b11111110, 
8'b00000010, 
8'b11111101, 
8'b00000001, 
8'b11111110, 
8'b00000000, 
8'b00000000, 
8'b11111100, 
8'b11111111, 
8'b00000000, 
8'b11111101, 
8'b00000000, 
8'b00000010, 
8'b11111110, 
8'b00000001, 
8'b11111111, 
8'b00000011, 
8'b11111010, 
8'b11111010, 
8'b00000001, 
8'b11111110, 
8'b00000000, 
8'b11111101, 
8'b11111111, 
8'b00000001, 
8'b00000000, 
8'b11111111, 
8'b00000000, 
8'b11111110, 
8'b00000010, 
8'b11111111, 
8'b11111110, 
8'b00000001, 
8'b11111111, 
8'b00000000, 
8'b00000001, 
8'b11111100, 
8'b11111110, 
8'b11111010, 
8'b00000001, 
8'b11111100, 
8'b00000001, 
8'b00000001, 
8'b11111111, 
8'b11111101, 
8'b11111110, 
8'b00000001, 
8'b11111111, 
8'b11111011, 
8'b00000011, 
8'b11111011, 
8'b11111101, 
8'b11111111, 
8'b00000000, 
8'b11111101, 
8'b11111110, 
8'b11111111, 
8'b11111111, 
8'b11111111, 
8'b11111111, 
8'b11111110, 
8'b00000011, 
8'b11111111, 
8'b00000000, 
8'b00000000, 
8'b11111111, 
8'b00000000, 
8'b00000000, 
8'b11111111, 
8'b11111111, 
8'b00000000, 
8'b00000000, 
8'b00000000, 
8'b00000001, 
8'b11111101, 
8'b00000011, 
8'b11111110, 
8'b00000000, 
8'b11111110, 
8'b00000001, 
8'b11111101, 
8'b11111101, 
8'b11111100, 
8'b11111111, 
8'b11111010, 
8'b11111111, 
8'b11111110, 
8'b11111101, 
8'b11111101, 
8'b11111110, 
8'b11111110, 
8'b00000010, 
8'b11111010, 
8'b00000100, 
8'b11111111, 
8'b11111101, 
8'b11111111, 
8'b11111100, 
8'b00000000, 
8'b00000001, 
8'b11111101, 
8'b00000000, 
8'b11111100, 
8'b00000010, 
8'b11111100, 
8'b00000000, 
8'b11111110, 
8'b11111111, 
8'b00000010, 
8'b00000010, 
8'b11111110, 
8'b00000010, 
8'b00000000, 
8'b00000000, 
8'b00000011, 
8'b00000001, 
8'b11111110, 
8'b11111110, 
8'b00000010, 
8'b00000010, 
8'b00000000, 
8'b00000001, 
8'b00000000, 
8'b00000000, 
8'b11111111, 
8'b00000010, 
8'b11111111, 
8'b00000000, 
8'b00000000, 
8'b00000100, 
8'b11111101, 
8'b11111110, 
8'b00000000, 
8'b00000010, 
8'b00000010, 
8'b11111101, 
8'b11111101, 
8'b00000000, 
8'b00000000, 
8'b00000000, 
8'b00000000, 
8'b00000001, 
8'b00000000, 
8'b00000010, 
8'b11111111, 
8'b00000000, 
8'b00000010, 
8'b11111111, 
8'b11111111, 
8'b00000000, 
8'b11111100, 
8'b00000000, 
8'b00000001, 
8'b11111101, 
8'b00000011, 
8'b11111111, 
8'b00000000, 
8'b11111111, 
8'b11111111, 
8'b11111111, 
8'b00000001, 
8'b00000011, 
8'b00000000, 
8'b00000001, 
8'b00000100, 
8'b11111100, 
8'b00000001, 
8'b00000010, 
8'b11111101, 
8'b00000000, 
8'b00000010, 
8'b00000000, 
8'b00000001, 
8'b11111111, 
8'b00000011, 
8'b00000001, 
8'b11111110, 
8'b11111100, 
8'b11111101, 
8'b00000000, 
8'b00000000, 
8'b11111111, 
8'b00000001, 
8'b00000001, 
8'b00000001, 
8'b11111100, 
8'b00000000, 
8'b00000001, 
8'b11111100, 
8'b11111110, 
8'b11111111, 
8'b00000011, 
8'b00000011, 
8'b11111111, 
8'b00000001, 
8'b11111100, 
8'b11111110, 
8'b11111110, 
8'b11111111, 
8'b00000000, 
8'b11111011, 
8'b00000001, 
8'b11111111, 
8'b11111111, 
8'b11111101, 
8'b00000000, 
8'b11111111, 
8'b00000100, 
8'b11111100, 
8'b00000001, 
8'b00000000, 
8'b11111110, 
8'b11111110, 
8'b00000000, 
8'b11111101, 
8'b11111110, 
8'b11111100, 
8'b11111111, 
8'b00000001, 
8'b00000011, 
8'b11111101, 
8'b11111111, 
8'b00000000, 
8'b00000010, 
8'b11111110, 
8'b11111111, 
8'b11111111, 
8'b00000010, 
8'b11111011, 
8'b00000010, 
8'b11111110, 
8'b11111011, 
8'b11111101, 
8'b00000100, 
8'b11111100, 
8'b11111111, 
8'b11111100, 
8'b00000001, 
8'b00000011, 
8'b00000011, 
8'b11111101, 
8'b00000000, 
8'b11111011, 
8'b00000001, 
8'b11111110, 
8'b00000010, 
8'b00000000, 
8'b00000001, 
8'b11111110, 
8'b11111110, 
8'b11111101, 
8'b00000000, 
8'b00000001, 
8'b00000011, 
8'b00000000, 
8'b11111110, 
8'b11111111, 
8'b11111100, 
8'b00000010, 
8'b00000001, 
8'b11111101, 
8'b11111111, 
8'b11111011, 
8'b00000010, 
8'b11111100, 
8'b00000011, 
8'b11111101, 
8'b00000000, 
8'b00000000, 
8'b00000010, 
8'b11111101, 
8'b11111101, 
8'b00000010, 
8'b11111110, 
8'b00000000, 
8'b11111101, 
8'b00000000, 
8'b11111110, 
8'b00000001, 
8'b11111110, 
8'b11111110, 
8'b11111110, 
8'b00000001, 
8'b11111110, 
8'b11111111, 
8'b00000001, 
8'b00000010, 
8'b11111100, 
8'b00000000, 
8'b00000000, 
8'b11111011, 
8'b11111111, 
8'b00000011, 
8'b00000001, 
8'b11111100, 
8'b00000001, 
8'b11111001, 
8'b11111100, 
8'b11111101, 
8'b00000000, 
8'b11111011, 
8'b11111110, 
8'b00000000, 
8'b11111110, 
8'b00000011, 
8'b00000000, 
8'b00000000, 
8'b00000000, 
8'b00000100, 
8'b11111101, 
8'b11111101, 
8'b00000000, 
8'b00000010, 
8'b00000010, 
8'b00000010, 
8'b11111110, 
8'b11111101, 
8'b00000000, 
8'b11111101, 
8'b00000000, 
8'b00000000, 
8'b00000000, 
8'b11111100, 
8'b11111100, 
8'b11111111, 
8'b11111111, 
8'b11111111, 
8'b11111100, 
8'b00000000, 
8'b11111110, 
8'b11111011, 
8'b11111101, 
8'b00000010, 
8'b11111100, 
8'b00000010, 
8'b00000100, 
8'b00000011, 
8'b11111111, 
8'b11111101, 
8'b00000001, 
8'b11111101, 
8'b11111110, 
8'b00000001, 
8'b11111111, 
8'b11111111, 
8'b11111111, 
8'b00000010
};
localparam logic signed [7:0] dlBiases [9:0] = {
8'b00000010, 
8'b11111111, 
8'b11111111, 
8'b11111111, 
8'b11111111, 
8'b11111111, 
8'b11111111, 
8'b00000001, 
8'b11111101, 
8'b11111111
};
localparam logic signed [7:0] convWeights [0:17] = {
8'b00000001, 
8'b00000111, 
8'b11111100, 
8'b00000001, 
8'b00000000, 
8'b00001000, 
8'b00000110, 
8'b00000011, 
8'b11111100, 
8'b00000101, 
8'b11111110, 
8'b00000011, 
8'b00000111, 
8'b00000010, 
8'b00000110, 
8'b11111111, 
8'b00000010, 
8'b00000001
};
localparam logic signed [7:0] convBiases [1:0] = {
8'b00000000, 
8'b00000000
};
endpackage