package data16_10;

//localparam logic [16:0] num = 17'b00000000001001000;
localparam logic signed [15:0] dlWeights [0:1279]= {
16'b0000000100000111, 
16'b0000000000001010, 
16'b1111111100111000, 
16'b0000000000000110, 
16'b1111111110111101, 
16'b0000000010001001, 
16'b0000000001000000, 
16'b1111111100110100, 
16'b0000000000101110, 
16'b0000000010101011, 
16'b0000000010101100, 
16'b1111111011110111, 
16'b1111111001111011, 
16'b1111111101010011, 
16'b0000000001100010, 
16'b1111111110000100, 
16'b1111111110110011, 
16'b1111111111100001, 
16'b1111111111001100, 
16'b1111111111111100, 
16'b0000000001111011, 
16'b1111111100001011, 
16'b0000000000110111, 
16'b0000000001010010, 
16'b1111111111011110, 
16'b0000000000000101, 
16'b1111111110111100, 
16'b0000000000100011, 
16'b0000000001000010, 
16'b0000000100000011, 
16'b0000001001001011, 
16'b1111111001001010, 
16'b1111111100000110, 
16'b1111111011010100, 
16'b1111111100010001, 
16'b0000000001111100, 
16'b1111111111100101, 
16'b0000000010100110, 
16'b1111111110110111, 
16'b0000000011010010, 
16'b0000000010011111, 
16'b1111111101110101, 
16'b1111111111101110, 
16'b1111111101010010, 
16'b0000000000000101, 
16'b1111111110011110, 
16'b0000000010110010, 
16'b1111111101100110, 
16'b1111111110001101, 
16'b0000000000001010, 
16'b0000000101110101, 
16'b1111111101101101, 
16'b1111111011111000, 
16'b1111111010101001, 
16'b1111111101011010, 
16'b0000000001100011, 
16'b1111111111101001, 
16'b0000000010000010, 
16'b0000000001000001, 
16'b0000000001101001, 
16'b0000000011111000, 
16'b1111111100110101, 
16'b0000000001000011, 
16'b0000000001000100, 
16'b1111111101010010, 
16'b0000000011101001, 
16'b0000000011011010, 
16'b0000000000000010, 
16'b0000000010110011, 
16'b1111111110101110, 
16'b0000000000000011, 
16'b0000000011010110, 
16'b1111111100011111, 
16'b1111111101100011, 
16'b1111111101011101, 
16'b0000000001100101, 
16'b1111111111010111, 
16'b0000000010110100, 
16'b1111111100010001, 
16'b1111111101000111, 
16'b1111111110110010, 
16'b1111111110010100, 
16'b1111111100011000, 
16'b0000000001101011, 
16'b1111111101110110, 
16'b0000000010001000, 
16'b0000000000000000, 
16'b1111111101010011, 
16'b1111111111000111, 
16'b1111111110001110, 
16'b0000000000100100, 
16'b0000000000010001, 
16'b1111111110010011, 
16'b0000000000011100, 
16'b1111111011100000, 
16'b1111111111001011, 
16'b1111111100001011, 
16'b0000000101000001, 
16'b1111111011110110, 
16'b1111111011001010, 
16'b0000000000010101, 
16'b0000000100110000, 
16'b0000000000000101, 
16'b0000000000100011, 
16'b1111111101100110, 
16'b1111111111100111, 
16'b1111111101001001, 
16'b1111111101010100, 
16'b0000000001101111, 
16'b1111111100111000, 
16'b0000000000011100, 
16'b0000000010101010, 
16'b0000000000100011, 
16'b0000000010000010, 
16'b1111111100000010, 
16'b1111111110011001, 
16'b1111111011110010, 
16'b0000000001110001, 
16'b1111111101010111, 
16'b0000000001000001, 
16'b1111111101000001, 
16'b1111111111000111, 
16'b0000000000010001, 
16'b0000000001001101, 
16'b1111111100001110, 
16'b1111111110111101, 
16'b1111111100010010, 
16'b1111111110011000, 
16'b0000000000000010, 
16'b0000000001010100, 
16'b1111111101011010, 
16'b1111111110111110, 
16'b1111111110010101, 
16'b0000000100011110, 
16'b1111111101001101, 
16'b1111111010111000, 
16'b1111111101101001, 
16'b0000000101000100, 
16'b1111111111001001, 
16'b0000000000110000, 
16'b1111111111110011, 
16'b1111111110101111, 
16'b0000000000001111, 
16'b0000000000110000, 
16'b0000000011001111, 
16'b1111111111010110, 
16'b1111111011110010, 
16'b0000000011010011, 
16'b1111111111001000, 
16'b0000000001000110, 
16'b0000000000010100, 
16'b0000000001010101, 
16'b0000000010010101, 
16'b1111111111110101, 
16'b0000000001010011, 
16'b1111111101101010, 
16'b1111110011111111, 
16'b0000000011001100, 
16'b1111111111010010, 
16'b0000000001100110, 
16'b0000000010100011, 
16'b1111111111000100, 
16'b1111111011110111, 
16'b0000000010111101, 
16'b0000000011011100, 
16'b1111111110010011, 
16'b0000000100000010, 
16'b1111111111000101, 
16'b0000000000101011, 
16'b1111111111101100, 
16'b0000000010010111, 
16'b1111111111110000, 
16'b1111111111000100, 
16'b1111111010100010, 
16'b0000000000010011, 
16'b0000000000111001, 
16'b1111111110101011, 
16'b1111111111100100, 
16'b1111111110001101, 
16'b0000000010010110, 
16'b0000000011110000, 
16'b1111111100010000, 
16'b1111111111101110, 
16'b1111111110100010, 
16'b0000000011110010, 
16'b1111111111110110, 
16'b0000000010001110, 
16'b1111111110001111, 
16'b0000000011001011, 
16'b0000000000000111, 
16'b0000000011110000, 
16'b1111111010011100, 
16'b1111111101101011, 
16'b1111111011110001, 
16'b1111111111111001, 
16'b0000000001011101, 
16'b0000000000101011, 
16'b0000000001101010, 
16'b0000000010011111, 
16'b1111111111010010, 
16'b0000000011010001, 
16'b1111111011110100, 
16'b1111111110010010, 
16'b1111111101110100, 
16'b1111111111111110, 
16'b0000000000001011, 
16'b0000000000000011, 
16'b1111111111011111, 
16'b0000000000010101, 
16'b1111111110011000, 
16'b1111111111000101, 
16'b1111111111010101, 
16'b1111111111010010, 
16'b1111111100101100, 
16'b1111111111110000, 
16'b0000000000011010, 
16'b0000000011010100, 
16'b1111111110100010, 
16'b0000000000001111, 
16'b0000000000101101, 
16'b1111111101110111, 
16'b1111111111001100, 
16'b1111111100111011, 
16'b0000000010111110, 
16'b1111111100110111, 
16'b0000000011110101, 
16'b1111111101001001, 
16'b0000000000010011, 
16'b1111111110101011, 
16'b1111111011101111, 
16'b0000000010100010, 
16'b0000000011101011, 
16'b1111111100111111, 
16'b0000000001000111, 
16'b1111111111101000, 
16'b0000000000001110, 
16'b1111111110010100, 
16'b0000000010100010, 
16'b0000000000111111, 
16'b0000000000110011, 
16'b0000000000000011, 
16'b1111111110010100, 
16'b0000000001010100, 
16'b0000000001111011, 
16'b0000000001010000, 
16'b1111111110101100, 
16'b1111111101010110, 
16'b1111111110111110, 
16'b0000000001111001, 
16'b1111111101101001, 
16'b0000000001001100, 
16'b0000000001000110, 
16'b1111111110110011, 
16'b1111111101111111, 
16'b1111111011110100, 
16'b1111111110010110, 
16'b0000000000001010, 
16'b0000000000000001, 
16'b1111111011001010, 
16'b1111111100101111, 
16'b1111111100000000, 
16'b0000000000101100, 
16'b0000000000011111, 
16'b0000000001011010, 
16'b1111111010101011, 
16'b0000000000010111, 
16'b0000000001110001, 
16'b1111111100101110, 
16'b0000000000001001, 
16'b1111111111100111, 
16'b0000000000011110, 
16'b0000000010111100, 
16'b0000000000110100, 
16'b0000000000011101, 
16'b1111111111011100, 
16'b1111111100110001, 
16'b1111111100011100, 
16'b0000000100001111, 
16'b1111111011100101, 
16'b0000000000010101, 
16'b1111111111110100, 
16'b0000000000001000, 
16'b0000000001011010, 
16'b1111111111001010, 
16'b0000000000100011, 
16'b1111111110010000, 
16'b0000000001101000, 
16'b1111111111111110, 
16'b0000000010010001, 
16'b0000000001011101, 
16'b1111111110010001, 
16'b0000000001110110, 
16'b0000000001110111, 
16'b0000000000000101, 
16'b0000000001011010, 
16'b1111111110011110, 
16'b1111111011001000, 
16'b1111111111101101, 
16'b1111111101010001, 
16'b1111111110111010, 
16'b0000000000100110, 
16'b0000000011001100, 
16'b0000000000110000, 
16'b0000000001011110, 
16'b1111111110111000, 
16'b0000000000101000, 
16'b0000000001010101, 
16'b1111111110111100, 
16'b0000000001100110, 
16'b0000000011001110, 
16'b0000000001111111, 
16'b0000000001001100, 
16'b1111111111011001, 
16'b0000000000110000, 
16'b0000000010010111, 
16'b0000000001010100, 
16'b1111111100001101, 
16'b0000000000010010, 
16'b1111111111010100, 
16'b1111111111111011, 
16'b0000000010000101, 
16'b1111111011101101, 
16'b1111111101110011, 
16'b0000000001101100, 
16'b0000000011011100, 
16'b0000000000010011, 
16'b0000000011011111, 
16'b1111111011111001, 
16'b0000000000001000, 
16'b0000000001111010, 
16'b0000000100011101, 
16'b1111111011110001, 
16'b1111111110101000, 
16'b1111111010111011, 
16'b1111111111000000, 
16'b0000000001100111, 
16'b1111111101111111, 
16'b0000000000101100, 
16'b1111111110100111, 
16'b1111111101101000, 
16'b0000000001111000, 
16'b1111111110101000, 
16'b1111111111001110, 
16'b1111111101000001, 
16'b0000000000100111, 
16'b1111111110111001, 
16'b0000000000111101, 
16'b1111111110010110, 
16'b0000000010100011, 
16'b1111111101110011, 
16'b0000000010100011, 
16'b1111111110110101, 
16'b1111111010011010, 
16'b0000000000110011, 
16'b0000000010011010, 
16'b0000000000001011, 
16'b0000000000011011, 
16'b0000000000100001, 
16'b0000000010100101, 
16'b1111111110011100, 
16'b0000000000101111, 
16'b1111111100000111, 
16'b0000000010000001, 
16'b0000000010010001, 
16'b0000000000010011, 
16'b1111111110111100, 
16'b0000000001010011, 
16'b1111111111000010, 
16'b0000000001000101, 
16'b0000000000100011, 
16'b0000000000000001, 
16'b0000000000011000, 
16'b1111111101100111, 
16'b0000000000110000, 
16'b1111111111010011, 
16'b0000000000100111, 
16'b0000000011010100, 
16'b0000000010001011, 
16'b1111111111101001, 
16'b1111111100110101, 
16'b0000000001110010, 
16'b1111111100010101, 
16'b1111111110111111, 
16'b1111111110011110, 
16'b1111111111111011, 
16'b0000000010101111, 
16'b1111111111001011, 
16'b0000000000000010, 
16'b0000000011111000, 
16'b1111111111010001, 
16'b1111111111010001, 
16'b1111111110111100, 
16'b1111111111101100, 
16'b0000000010000100, 
16'b1111111101001000, 
16'b1111111110100111, 
16'b1111111110101010, 
16'b1111111100111010, 
16'b1111111101111000, 
16'b1111111011110100, 
16'b1111111110010110, 
16'b1111111110011100, 
16'b1111111011111111, 
16'b0000000011000110, 
16'b1111111100111111, 
16'b0000000001000110, 
16'b1111111101010111, 
16'b1111111101011001, 
16'b0000000001111011, 
16'b0000000000000011, 
16'b1111111101001010, 
16'b0000000000101110, 
16'b1111111100101110, 
16'b0000000010100100, 
16'b0000000001001000, 
16'b1111111110110100, 
16'b1111111101111011, 
16'b1111111110000011, 
16'b0000000001100111, 
16'b1111111101000000, 
16'b0000000000001010, 
16'b0000000010100100, 
16'b0000000001011000, 
16'b0000000001101101, 
16'b1111111101001100, 
16'b0000000011001111, 
16'b0000000010011101, 
16'b0000000000011001, 
16'b0000000011101000, 
16'b0000000000011101, 
16'b1111111011100111, 
16'b0000000011011000, 
16'b0000000001010011, 
16'b0000000010110011, 
16'b1111111100011100, 
16'b1111111111010011, 
16'b0000000000111001, 
16'b1111111101001110, 
16'b1111111101100100, 
16'b1111111101101110, 
16'b1111111110010111, 
16'b0000000011101010, 
16'b0000000000001101, 
16'b0000000001101000, 
16'b0000000000001100, 
16'b0000000011000010, 
16'b0000000010111000, 
16'b1111111100001111, 
16'b1111111101011000, 
16'b0000000010001101, 
16'b1111111101111011, 
16'b1111111111011000, 
16'b1111111111011000, 
16'b0000000010000011, 
16'b0000000000110001, 
16'b1111111111110111, 
16'b1111111101010101, 
16'b0000000010011110, 
16'b1111111111001010, 
16'b0000000010101110, 
16'b0000000000111101, 
16'b0000000001010101, 
16'b1111111110111110, 
16'b0000000000010001, 
16'b0000000010101110, 
16'b1111111111011101, 
16'b1111111111110100, 
16'b1111111111101000, 
16'b1111111101100111, 
16'b0000000100000001, 
16'b0000000000100110, 
16'b1111111110000101, 
16'b1111111111101010, 
16'b0000000000111000, 
16'b1111111111010011, 
16'b1111111111010001, 
16'b0000000000100100, 
16'b0000000011001011, 
16'b0000000001110001, 
16'b0000000010110110, 
16'b0000000000111111, 
16'b1111111101101000, 
16'b0000000000101000, 
16'b1111111101101000, 
16'b1111111110101010, 
16'b1111111110000100, 
16'b0000000000000001, 
16'b0000000000010110, 
16'b0000000001010111, 
16'b0000000000110011, 
16'b0000000001000001, 
16'b1111111011001110, 
16'b1111111101100000, 
16'b1111111111100001, 
16'b0000000000011100, 
16'b0000000011110110, 
16'b0000000011110001, 
16'b1111111011110011, 
16'b1111111111011111, 
16'b0000000010000100, 
16'b0000000011010110, 
16'b1111111011110011, 
16'b1111111101101001, 
16'b0000000000011100, 
16'b0000000010010110, 
16'b1111111110100011, 
16'b1111111110111011, 
16'b1111111111001001, 
16'b1111111111110101, 
16'b0000000011010110, 
16'b0000000010101001, 
16'b1111111111101101, 
16'b1111111110110110, 
16'b0000000010010110, 
16'b0000000001001000, 
16'b0000000010001010, 
16'b1111111111100111, 
16'b1111111110000111, 
16'b1111111111000110, 
16'b1111111111100100, 
16'b1111111100101000, 
16'b0000000000101101, 
16'b1111111100110000, 
16'b0000000001100111, 
16'b1111111111100001, 
16'b1111111111100101, 
16'b0000000010000011, 
16'b0000000000010011, 
16'b1111111111101011, 
16'b0000000001010110, 
16'b0000000001000011, 
16'b0000000000110111, 
16'b0000000000011011, 
16'b0000000001100000, 
16'b1111111101111101, 
16'b0000000100000010, 
16'b0000000001111110, 
16'b1111111011101001, 
16'b0000000000010010, 
16'b1111111100100001, 
16'b1111111100011000, 
16'b1111111011010111, 
16'b1111111111001010, 
16'b1111111110101011, 
16'b1111111110000011, 
16'b0000000001011011, 
16'b0000000000010000, 
16'b1111111100111110, 
16'b0000000000101001, 
16'b1111111110000110, 
16'b1111111110010000, 
16'b1111111110100000, 
16'b1111111110111101, 
16'b1111111110011000, 
16'b0000000000010001, 
16'b1111111111001001, 
16'b0000000010010110, 
16'b1111111110000001, 
16'b0000000000110110, 
16'b0000000000011001, 
16'b0000000001011001, 
16'b0000000011011001, 
16'b0000000000000001, 
16'b1111111101110101, 
16'b1111111110100000, 
16'b0000000001110010, 
16'b0000000010001110, 
16'b1111111010111101, 
16'b0000000001001101, 
16'b0000000000010011, 
16'b1111111011101010, 
16'b0000000010110101, 
16'b1111111110110001, 
16'b0000000000000100, 
16'b1111111101101110, 
16'b0000000010110000, 
16'b0000000001111100, 
16'b1111111010011010, 
16'b0000000010001110, 
16'b0000000001011111, 
16'b0000000001011001, 
16'b0000000100101001, 
16'b0000000001010011, 
16'b0000000010100010, 
16'b1111111101100011, 
16'b0000000000100100, 
16'b1111111111000100, 
16'b0000000001000100, 
16'b0000000011101100, 
16'b0000000001110110, 
16'b1111111010111010, 
16'b0000000010100110, 
16'b1111111110110110, 
16'b0000000000101101, 
16'b1111111101111101, 
16'b1111111101001001, 
16'b0000000000100011, 
16'b0000000001111000, 
16'b0000000000111101, 
16'b1111111111000110, 
16'b1111111011011000, 
16'b0000000001001010, 
16'b0000000000011011, 
16'b0000000010010100, 
16'b0000000000000110, 
16'b0000000000100010, 
16'b0000000010011101, 
16'b0000000010001000, 
16'b1111111110110110, 
16'b0000000001101110, 
16'b1111111101111101, 
16'b1111111101111110, 
16'b1111111110101000, 
16'b0000000010110010, 
16'b1111111110000111, 
16'b1111111101001111, 
16'b0000000000011101, 
16'b0000000001101111, 
16'b0000000010001001, 
16'b1111111110011101, 
16'b1111111011101110, 
16'b1111111011100111, 
16'b0000000001111010, 
16'b0000000000001111, 
16'b0000000010101110, 
16'b0000000010001101, 
16'b0000000001110111, 
16'b0000000010111000, 
16'b1111111110100111, 
16'b1111111111110000, 
16'b0000000000101101, 
16'b0000000001001010, 
16'b0000000010011100, 
16'b0000000010101110, 
16'b0000000011010000, 
16'b1111111101111001, 
16'b0000000000000001, 
16'b0000000011010100, 
16'b0000000010011011, 
16'b0000000010010001, 
16'b1111111111110011, 
16'b1111111101011111, 
16'b1111111111010100, 
16'b1111111111011010, 
16'b1111111101111000, 
16'b1111111100000100, 
16'b0000000010000111, 
16'b0000000001111000, 
16'b0000000010100001, 
16'b0000000000000010, 
16'b1111111110011110, 
16'b1111111111010111, 
16'b1111111110000110, 
16'b0000000000011110, 
16'b0000000000000010, 
16'b0000000010111101, 
16'b0000000001010011, 
16'b1111111011100010, 
16'b1111111101101110, 
16'b1111111101001011, 
16'b1111111111111001, 
16'b1111111100011000, 
16'b1111111111001111, 
16'b1111111110110100, 
16'b0000000000110111, 
16'b0000000000001001, 
16'b0000000000100011, 
16'b1111111011001101, 
16'b1111111111110100, 
16'b0000000010001010, 
16'b0000000011011000, 
16'b1111111111101010, 
16'b1111111100001111, 
16'b0000000001111001, 
16'b1111111111000110, 
16'b0000000010110101, 
16'b1111111111111010, 
16'b1111111011011111, 
16'b1111111110100001, 
16'b0000000000010110, 
16'b1111111100010011, 
16'b1111111111101010, 
16'b0000000010110100, 
16'b1111111110110100, 
16'b1111111111110101, 
16'b0000000010101111, 
16'b0000000000111011, 
16'b1111111110110111, 
16'b0000000010111000, 
16'b1111111110111000, 
16'b0000000001001100, 
16'b0000000000001101, 
16'b1111111100111010, 
16'b0000000010100001, 
16'b1111111110011011, 
16'b0000000000001001, 
16'b0000000000010100, 
16'b1111111110100111, 
16'b1111111111001100, 
16'b0000000001110001, 
16'b0000000000000010, 
16'b0000000000101101, 
16'b0000000001001101, 
16'b1111111110001110, 
16'b0000000000111010, 
16'b1111111101010110, 
16'b1111111111111011, 
16'b1111111110011011, 
16'b1111111110010100, 
16'b1111111101100100, 
16'b0000000000011000, 
16'b0000000001010100, 
16'b0000000000101111, 
16'b1111111110110000, 
16'b1111111101101010, 
16'b0000000010101001, 
16'b1111111110011111, 
16'b0000000000000001, 
16'b0000000011001111, 
16'b0000000000000100, 
16'b1111111100110010, 
16'b0000000010001101, 
16'b1111111101110011, 
16'b0000000001011101, 
16'b0000000000111111, 
16'b0000000001000001, 
16'b0000000010000111, 
16'b1111111101100001, 
16'b0000000000110010, 
16'b1111111110011000, 
16'b1111111101000101, 
16'b0000000001101110, 
16'b1111111100111010, 
16'b0000000010110101, 
16'b0000000000100010, 
16'b1111111110111000, 
16'b1111111100110010, 
16'b1111111110100111, 
16'b0000000010101001, 
16'b1111111110000011, 
16'b0000000000001010, 
16'b1111111110101001, 
16'b0000000011000000, 
16'b1111111111011110, 
16'b0000000000010011, 
16'b0000000001100001, 
16'b1111111110011010, 
16'b1111111110001100, 
16'b0000000000110000, 
16'b0000000000011001, 
16'b1111111100010100, 
16'b0000000011011010, 
16'b1111111111010010, 
16'b0000000011001010, 
16'b0000000001110001, 
16'b0000000001100100, 
16'b1111111101110000, 
16'b1111111111010000, 
16'b1111111111010000, 
16'b1111111110111000, 
16'b1111111111101011, 
16'b0000000001110001, 
16'b1111111110000011, 
16'b0000000001100110, 
16'b0000000000010111, 
16'b0000000000100010, 
16'b0000000001101001, 
16'b0000000010100001, 
16'b0000000001010101, 
16'b1111111110001000, 
16'b0000000000111010, 
16'b1111111100001111, 
16'b0000000001000100, 
16'b1111111110110100, 
16'b0000000001100010, 
16'b1111111110100100, 
16'b1111111110010011, 
16'b0000000001010101, 
16'b1111111101100011, 
16'b1111111110011111, 
16'b1111111101010011, 
16'b0000000000011101, 
16'b1111111110001101, 
16'b0000000011100110, 
16'b1111111111101001, 
16'b1111111110001000, 
16'b1111111111111100, 
16'b0000000001010010, 
16'b0000000001010000, 
16'b0000000010101111, 
16'b1111111110101111, 
16'b1111111101000000, 
16'b0000000000001101, 
16'b1111111101111011, 
16'b1111111110101110, 
16'b1111111100100000, 
16'b0000000001101100, 
16'b0000000100001101, 
16'b0000000001100111, 
16'b0000000010100111, 
16'b1111111111111001, 
16'b1111111110001100, 
16'b0000000010010000, 
16'b1111111111000011, 
16'b0000000010100011, 
16'b1111111110110011, 
16'b0000000000101110, 
16'b1111111101000110, 
16'b0000000100011000, 
16'b0000000011110010, 
16'b1111111110010011, 
16'b1111111010111001, 
16'b0000000000010111, 
16'b1111111101100011, 
16'b0000000100000011, 
16'b1111111111100000, 
16'b1111111110011011, 
16'b0000000000011010, 
16'b1111111110001100, 
16'b1111111110010101, 
16'b1111111110111011, 
16'b1111111011001111, 
16'b0000000000011110, 
16'b1111111011010100, 
16'b1111111110101010, 
16'b0000000000011011, 
16'b0000000001011101, 
16'b1111111110001111, 
16'b1111111111101110, 
16'b0000000000101000, 
16'b1111111110110110, 
16'b1111111010101000, 
16'b1111111110110101, 
16'b0000000000110101, 
16'b0000000000100101, 
16'b0000000001001010, 
16'b0000000001010001, 
16'b1111111011101110, 
16'b1111111110100000, 
16'b0000000010110001, 
16'b1111111100111001, 
16'b1111111110111000, 
16'b0000000011101110, 
16'b1111111110011000, 
16'b0000000000000110, 
16'b1111111110011100, 
16'b0000000000100001, 
16'b1111111111010111, 
16'b1111111110111001, 
16'b0000000010111110, 
16'b1111111100111111, 
16'b1111111110111001, 
16'b0000000010010010, 
16'b0000000010111010, 
16'b1111111111001010, 
16'b0000000001000010, 
16'b1111111111011000, 
16'b1111111011101000, 
16'b1111111110111100, 
16'b0000000000100100, 
16'b1111111110011100, 
16'b1111111111111000, 
16'b1111111111000000, 
16'b1111111110011100, 
16'b0000000010011010, 
16'b1111111110011101, 
16'b1111111110000000, 
16'b0000000000001100, 
16'b1111111111000000, 
16'b0000000001010001, 
16'b1111111101011000, 
16'b0000000010100000, 
16'b0000000001111111, 
16'b0000000000001011, 
16'b1111111111111010, 
16'b1111111101110001, 
16'b1111111101010110, 
16'b1111111110001100, 
16'b1111111110110110, 
16'b1111111111011110, 
16'b0000000000101000, 
16'b0000000011110011, 
16'b1111111110111010, 
16'b1111111100011101, 
16'b0000000011101011, 
16'b1111111110001101, 
16'b1111111111100100, 
16'b0000000000100010, 
16'b0000000001101011, 
16'b1111111101111101, 
16'b1111111110001000, 
16'b1111111111001100, 
16'b0000000001110111, 
16'b1111111110011101, 
16'b0000000001100101, 
16'b0000000001110101, 
16'b1111111101001100, 
16'b0000000000000111, 
16'b0000000000000011, 
16'b1111111111001100, 
16'b1111111110110010, 
16'b0000000000010110, 
16'b1111111111001110, 
16'b0000000000111001, 
16'b0000000000110110, 
16'b1111111101010010, 
16'b1111111110001001, 
16'b0000000000011101, 
16'b0000000001111000, 
16'b1111111100100001, 
16'b1111111011100111, 
16'b1111111110011100, 
16'b1111111111010011, 
16'b1111111111011110, 
16'b1111111111101101, 
16'b1111111101101101, 
16'b0000000001010110, 
16'b0000000001011110, 
16'b1111111110011101, 
16'b0000000001101101, 
16'b1111111111110001, 
16'b1111111110111010, 
16'b0000000010110001, 
16'b1111111110000111, 
16'b1111111111011011, 
16'b1111111110000110, 
16'b0000000000110010, 
16'b0000000010010001, 
16'b1111111111111000, 
16'b0000000001011011, 
16'b1111111011011100, 
16'b0000000000011011, 
16'b1111111110010111, 
16'b1111111110101100, 
16'b0000000010011010, 
16'b1111111101000111, 
16'b0000000001010100, 
16'b1111111110101111, 
16'b0000000000000100, 
16'b0000000000000100, 
16'b1111111100110010, 
16'b1111111111110011, 
16'b0000000000011110, 
16'b1111111101101101, 
16'b0000000000100000, 
16'b0000000010100000, 
16'b1111111110010001, 
16'b0000000001111001, 
16'b1111111111000111, 
16'b0000000011011110, 
16'b1111111010111110, 
16'b1111111010110001, 
16'b0000000001100011, 
16'b1111111110100100, 
16'b0000000000101010, 
16'b1111111101110111, 
16'b1111111111010111, 
16'b0000000001110110, 
16'b0000000000100010, 
16'b1111111111111000, 
16'b0000000000100000, 
16'b1111111110010010, 
16'b0000000010001011, 
16'b1111111111111011, 
16'b1111111110011101, 
16'b0000000001010001, 
16'b1111111111100010, 
16'b0000000000001110, 
16'b0000000001111101, 
16'b1111111100100111, 
16'b1111111110000001, 
16'b1111111010111101, 
16'b0000000001000000, 
16'b1111111100100101, 
16'b0000000001100000, 
16'b0000000001001111, 
16'b1111111111111111, 
16'b1111111101111110, 
16'b1111111110010111, 
16'b0000000001110011, 
16'b1111111111101001, 
16'b1111111011111100, 
16'b0000000011001011, 
16'b1111111011100010, 
16'b1111111101100110, 
16'b1111111111100001, 
16'b0000000000000001, 
16'b1111111101001001, 
16'b1111111110101101, 
16'b1111111111111100, 
16'b1111111111101101, 
16'b1111111111010000, 
16'b1111111111110101, 
16'b1111111110001011, 
16'b0000000011100011, 
16'b1111111111000100, 
16'b0000000000011100, 
16'b0000000000011101, 
16'b1111111111011000, 
16'b0000000000101001, 
16'b0000000000010111, 
16'b1111111111001111, 
16'b1111111111010011, 
16'b0000000000110110, 
16'b0000000000011010, 
16'b0000000000101100, 
16'b0000000001010110, 
16'b1111111101101000, 
16'b0000000011111001, 
16'b1111111110100001, 
16'b0000000000100001, 
16'b1111111110101000, 
16'b0000000001010011, 
16'b1111111101001110, 
16'b1111111101110011, 
16'b1111111100011101, 
16'b1111111111010100, 
16'b1111111010110010, 
16'b1111111111110110, 
16'b1111111110001111, 
16'b1111111101001000, 
16'b1111111101111000, 
16'b1111111110111110, 
16'b1111111110001000, 
16'b0000000010101000, 
16'b1111111010111101, 
16'b0000000100001000, 
16'b1111111111010111, 
16'b1111111101111011, 
16'b1111111111010101, 
16'b1111111100111011, 
16'b0000000000100100, 
16'b0000000001011000, 
16'b1111111101010110, 
16'b0000000000101110, 
16'b1111111100010010, 
16'b0000000010000100, 
16'b1111111100111111, 
16'b0000000000101111, 
16'b1111111110100010, 
16'b1111111111000011, 
16'b0000000010110010, 
16'b0000000010010010, 
16'b1111111110011000, 
16'b0000000010001111, 
16'b0000000000111000, 
16'b0000000000100110, 
16'b0000000011011010, 
16'b0000000001111101, 
16'b1111111110010000, 
16'b1111111110000001, 
16'b0000000010111000, 
16'b0000000010101011, 
16'b0000000000001110, 
16'b0000000001100001, 
16'b0000000000101111, 
16'b0000000000101101, 
16'b1111111111011000, 
16'b0000000010011110, 
16'b1111111111100001, 
16'b0000000000000011, 
16'b0000000000111101, 
16'b0000000100110010, 
16'b1111111101010110, 
16'b1111111110111011, 
16'b0000000000000111, 
16'b0000000010000000, 
16'b0000000010011111, 
16'b1111111101100011, 
16'b1111111101011000, 
16'b0000000000010100, 
16'b0000000000111001, 
16'b0000000000010100, 
16'b0000000000100001, 
16'b0000000001001000, 
16'b0000000000111010, 
16'b0000000010000100, 
16'b1111111111111001, 
16'b0000000000010110, 
16'b0000000010010000, 
16'b1111111111110110, 
16'b1111111111010001, 
16'b0000000000100001, 
16'b1111111100110011, 
16'b0000000000011000, 
16'b0000000001011001, 
16'b1111111101011101, 
16'b0000000011111011, 
16'b1111111111110001, 
16'b0000000000111110, 
16'b1111111111110101, 
16'b1111111111011011, 
16'b1111111111010010, 
16'b0000000001110111, 
16'b0000000011111100, 
16'b0000000000000000, 
16'b0000000001100001, 
16'b0000000100000010, 
16'b1111111100111100, 
16'b0000000001111000, 
16'b0000000010000011, 
16'b1111111101111011, 
16'b0000000000011111, 
16'b0000000010011101, 
16'b0000000000001111, 
16'b0000000001110100, 
16'b1111111111101110, 
16'b0000000011011100, 
16'b0000000001011110, 
16'b1111111110100011, 
16'b1111111100001110, 
16'b1111111101101110, 
16'b0000000000110010, 
16'b0000000000001110, 
16'b1111111111100001, 
16'b0000000001000111, 
16'b0000000001011010, 
16'b0000000001010100, 
16'b1111111100011001, 
16'b0000000000101111, 
16'b0000000001101001, 
16'b1111111100110110, 
16'b1111111110010111, 
16'b1111111111011101, 
16'b0000000011001001, 
16'b0000000011010101, 
16'b1111111111111100, 
16'b0000000001110101, 
16'b1111111100110101, 
16'b1111111110110101, 
16'b1111111110111100, 
16'b1111111111100101, 
16'b0000000000010010, 
16'b1111111011110000, 
16'b0000000001110110, 
16'b1111111111001011, 
16'b1111111111001000, 
16'b1111111101010000, 
16'b0000000000011101, 
16'b1111111111110111, 
16'b0000000100101111, 
16'b1111111100010111, 
16'b0000000001000000, 
16'b0000000000000111, 
16'b1111111110000101, 
16'b1111111110110010, 
16'b0000000000101001, 
16'b1111111101010110, 
16'b1111111110011101, 
16'b1111111100011110, 
16'b1111111111000110, 
16'b0000000001101110, 
16'b0000000011001100, 
16'b1111111101111011, 
16'b1111111111001100, 
16'b0000000000100110, 
16'b0000000010100101, 
16'b1111111110111101, 
16'b1111111111111100, 
16'b1111111111101010, 
16'b0000000010110001, 
16'b1111111011101110, 
16'b0000000010101011, 
16'b1111111110010000, 
16'b1111111011111001, 
16'b1111111101111000, 
16'b0000000100001010, 
16'b1111111100101110, 
16'b1111111111000100, 
16'b1111111100000010, 
16'b0000000001100011, 
16'b0000000011100001, 
16'b0000000011101100, 
16'b1111111101111100, 
16'b0000000000001100, 
16'b1111111011110010, 
16'b0000000001101101, 
16'b1111111110000100, 
16'b0000000010010111, 
16'b0000000000000101, 
16'b0000000001010000, 
16'b1111111110000010, 
16'b1111111110011011, 
16'b1111111101110111, 
16'b0000000000110011, 
16'b0000000001000110, 
16'b0000000011011111, 
16'b0000000000100010, 
16'b1111111110000101, 
16'b1111111111000011, 
16'b1111111100100100, 
16'b0000000010101010, 
16'b0000000001110110, 
16'b1111111101000100, 
16'b1111111111001110, 
16'b1111111011110011, 
16'b0000000010101011, 
16'b1111111100110010, 
16'b0000000011010001, 
16'b1111111101111110, 
16'b0000000000110001, 
16'b0000000000011011, 
16'b0000000010100001, 
16'b1111111101101111, 
16'b1111111101011111, 
16'b0000000010110100, 
16'b1111111110011011, 
16'b0000000000010100, 
16'b1111111101010100, 
16'b0000000000001100, 
16'b1111111110100001, 
16'b0000000001110101, 
16'b1111111110110101, 
16'b1111111110011010, 
16'b1111111110100001, 
16'b0000000001100100, 
16'b1111111110110010, 
16'b1111111111010101, 
16'b0000000001010001, 
16'b0000000010011011, 
16'b1111111100001011, 
16'b0000000000010010, 
16'b0000000000011011, 
16'b1111111011111001, 
16'b1111111111011001, 
16'b0000000011000101, 
16'b0000000001110100, 
16'b1111111100011101, 
16'b0000000001111011, 
16'b1111111001000100, 
16'b1111111100101111, 
16'b1111111101001010, 
16'b0000000000010000, 
16'b1111111011101010, 
16'b1111111110111001, 
16'b0000000000010010, 
16'b1111111110100000, 
16'b0000000011111111, 
16'b0000000000100000, 
16'b0000000000001010, 
16'b0000000000000000, 
16'b0000000100101100, 
16'b1111111101001110, 
16'b1111111101011111, 
16'b0000000000101110, 
16'b0000000010101000, 
16'b0000000010000001, 
16'b0000000010000011, 
16'b1111111110001010, 
16'b1111111101011110, 
16'b0000000000011110, 
16'b1111111101110101, 
16'b0000000000101011, 
16'b0000000000111110, 
16'b0000000000010100, 
16'b1111111100010111, 
16'b1111111100010101, 
16'b1111111111100100, 
16'b1111111111000111, 
16'b1111111111011011, 
16'b1111111100000101, 
16'b0000000000101011, 
16'b1111111110101001, 
16'b1111111011010101, 
16'b1111111101111010, 
16'b0000000010101110, 
16'b1111111100111101, 
16'b0000000010010011, 
16'b0000000100000010, 
16'b0000000011111100, 
16'b1111111111111000, 
16'b1111111101010111, 
16'b0000000001101111, 
16'b1111111101011000, 
16'b1111111110111000, 
16'b0000000001100111, 
16'b1111111111100100, 
16'b1111111111011111, 
16'b1111111111011011, 
16'b0000000010000011
};

localparam logic signed [15:0] dlBiases [9:0] = {
16'h00aa,
16'hfffe,
16'hfffe,
16'hffc4,
16'hffc1,
16'hffeb,
16'hffe9,
16'h004e,
16'hff47,
16'hffeb
};

localparam logic signed [15:0] convWeights [0:17] = {
16'b0000000001110010,
16'b0000000111101100,
16'b1111111100001011,
16'b0000000001011111,
16'b0000000000001110,
16'b0000001000001101,
16'b0000000110011111,
16'b0000000011001100,
16'b1111111100010110,
16'b0000000101100100,
16'b1111111110100111,
16'b0000000011010111,
16'b0000000111111101,
16'b0000000010100011,
16'b0000000110001000,
16'b1111111111110100,
16'b0000000010111010,
16'b0000000001110100 
};
localparam logic signed [15:0] convBiases  [1:0] = {
16'b0000000000000000,
16'b0000000000000000
};
endpackage