package data18_9;
localparam logic signed [17:0] dlWeights [0:1279] = {
18'b000000000010000011, 
18'b000000000000000101, 
18'b111111111110011100, 
18'b000000000000000011, 
18'b111111111111011110, 
18'b000000000001000100, 
18'b000000000000100000, 
18'b111111111110011010, 
18'b000000000000010111, 
18'b000000000001010101, 
18'b000000000001010110, 
18'b111111111101111011, 
18'b111111111100111101, 
18'b111111111110101001, 
18'b000000000000110001, 
18'b111111111111000010, 
18'b111111111111011001, 
18'b111111111111110000, 
18'b111111111111100110, 
18'b111111111111111110, 
18'b000000000000111101, 
18'b111111111110000101, 
18'b000000000000011011, 
18'b000000000000101001, 
18'b111111111111101111, 
18'b000000000000000010, 
18'b111111111111011110, 
18'b000000000000010001, 
18'b000000000000100001, 
18'b000000000010000001, 
18'b000000000100100101, 
18'b111111111100100101, 
18'b111111111110000011, 
18'b111111111101101010, 
18'b111111111110001000, 
18'b000000000000111110, 
18'b111111111111110010, 
18'b000000000001010011, 
18'b111111111111011011, 
18'b000000000001101001, 
18'b000000000001001111, 
18'b111111111110111010, 
18'b111111111111110111, 
18'b111111111110101001, 
18'b000000000000000010, 
18'b111111111111001111, 
18'b000000000001011001, 
18'b111111111110110011, 
18'b111111111111000110, 
18'b000000000000000101, 
18'b000000000010111010, 
18'b111111111110110110, 
18'b111111111101111100, 
18'b111111111101010100, 
18'b111111111110101101, 
18'b000000000000110001, 
18'b111111111111110100, 
18'b000000000001000001, 
18'b000000000000100000, 
18'b000000000000110100, 
18'b000000000001111100, 
18'b111111111110011010, 
18'b000000000000100001, 
18'b000000000000100010, 
18'b111111111110101001, 
18'b000000000001110100, 
18'b000000000001101101, 
18'b000000000000000001, 
18'b000000000001011001, 
18'b111111111111010111, 
18'b000000000000000001, 
18'b000000000001101011, 
18'b111111111110001111, 
18'b111111111110110001, 
18'b111111111110101110, 
18'b000000000000110010, 
18'b111111111111101011, 
18'b000000000001011010, 
18'b111111111110001000, 
18'b111111111110100011, 
18'b111111111111011001, 
18'b111111111111001010, 
18'b111111111110001100, 
18'b000000000000110101, 
18'b111111111110111011, 
18'b000000000001000100, 
18'b000000000000000000, 
18'b111111111110101001, 
18'b111111111111100011, 
18'b111111111111000111, 
18'b000000000000010010, 
18'b000000000000001000, 
18'b111111111111001001, 
18'b000000000000001110, 
18'b111111111101110000, 
18'b111111111111100101, 
18'b111111111110000101, 
18'b000000000010100000, 
18'b111111111101111011, 
18'b111111111101100101, 
18'b000000000000001010, 
18'b000000000010011000, 
18'b000000000000000010, 
18'b000000000000010001, 
18'b111111111110110011, 
18'b111111111111110011, 
18'b111111111110100100, 
18'b111111111110101010, 
18'b000000000000110111, 
18'b111111111110011100, 
18'b000000000000001110, 
18'b000000000001010101, 
18'b000000000000010001, 
18'b000000000001000001, 
18'b111111111110000001, 
18'b111111111111001100, 
18'b111111111101111001, 
18'b000000000000111000, 
18'b111111111110101011, 
18'b000000000000100000, 
18'b111111111110100000, 
18'b111111111111100011, 
18'b000000000000001000, 
18'b000000000000100110, 
18'b111111111110000111, 
18'b111111111111011110, 
18'b111111111110001001, 
18'b111111111111001100, 
18'b000000000000000001, 
18'b000000000000101010, 
18'b111111111110101101, 
18'b111111111111011111, 
18'b111111111111001010, 
18'b000000000010001111, 
18'b111111111110100110, 
18'b111111111101011100, 
18'b111111111110110100, 
18'b000000000010100010, 
18'b111111111111100100, 
18'b000000000000011000, 
18'b111111111111111001, 
18'b111111111111010111, 
18'b000000000000000111, 
18'b000000000000011000, 
18'b000000000001100111, 
18'b111111111111101011, 
18'b111111111101111001, 
18'b000000000001101001, 
18'b111111111111100100, 
18'b000000000000100011, 
18'b000000000000001010, 
18'b000000000000101010, 
18'b000000000001001010, 
18'b111111111111111010, 
18'b000000000000101001, 
18'b111111111110110101, 
18'b111111111001111111, 
18'b000000000001100110, 
18'b111111111111101001, 
18'b000000000000110011, 
18'b000000000001010001, 
18'b111111111111100010, 
18'b111111111101111011, 
18'b000000000001011110, 
18'b000000000001101110, 
18'b111111111111001001, 
18'b000000000010000001, 
18'b111111111111100010, 
18'b000000000000010101, 
18'b111111111111110110, 
18'b000000000001001011, 
18'b111111111111111000, 
18'b111111111111100010, 
18'b111111111101010001, 
18'b000000000000001001, 
18'b000000000000011100, 
18'b111111111111010101, 
18'b111111111111110010, 
18'b111111111111000110, 
18'b000000000001001011, 
18'b000000000001111000, 
18'b111111111110001000, 
18'b111111111111110111, 
18'b111111111111010001, 
18'b000000000001111001, 
18'b111111111111111011, 
18'b000000000001000111, 
18'b111111111111000111, 
18'b000000000001100101, 
18'b000000000000000011, 
18'b000000000001111000, 
18'b111111111101001110, 
18'b111111111110110101, 
18'b111111111101111000, 
18'b111111111111111100, 
18'b000000000000101110, 
18'b000000000000010101, 
18'b000000000000110101, 
18'b000000000001001111, 
18'b111111111111101001, 
18'b000000000001101000, 
18'b111111111101111010, 
18'b111111111111001001, 
18'b111111111110111010, 
18'b111111111111111111, 
18'b000000000000000101, 
18'b000000000000000001, 
18'b111111111111101111, 
18'b000000000000001010, 
18'b111111111111001100, 
18'b111111111111100010, 
18'b111111111111101010, 
18'b111111111111101001, 
18'b111111111110010110, 
18'b111111111111111000, 
18'b000000000000001101, 
18'b000000000001101010, 
18'b111111111111010001, 
18'b000000000000000111, 
18'b000000000000010110, 
18'b111111111110111011, 
18'b111111111111100110, 
18'b111111111110011101, 
18'b000000000001011111, 
18'b111111111110011011, 
18'b000000000001111010, 
18'b111111111110100100, 
18'b000000000000001001, 
18'b111111111111010101, 
18'b111111111101110111, 
18'b000000000001010001, 
18'b000000000001110101, 
18'b111111111110011111, 
18'b000000000000100011, 
18'b111111111111110100, 
18'b000000000000000111, 
18'b111111111111001010, 
18'b000000000001010001, 
18'b000000000000011111, 
18'b000000000000011001, 
18'b000000000000000001, 
18'b111111111111001010, 
18'b000000000000101010, 
18'b000000000000111101, 
18'b000000000000101000, 
18'b111111111111010110, 
18'b111111111110101011, 
18'b111111111111011111, 
18'b000000000000111100, 
18'b111111111110110100, 
18'b000000000000100110, 
18'b000000000000100011, 
18'b111111111111011001, 
18'b111111111110111111, 
18'b111111111101111010, 
18'b111111111111001011, 
18'b000000000000000101, 
18'b000000000000000000, 
18'b111111111101100101, 
18'b111111111110010111, 
18'b111111111110000000, 
18'b000000000000010110, 
18'b000000000000001111, 
18'b000000000000101101, 
18'b111111111101010101, 
18'b000000000000001011, 
18'b000000000000111000, 
18'b111111111110010111, 
18'b000000000000000100, 
18'b111111111111110011, 
18'b000000000000001111, 
18'b000000000001011110, 
18'b000000000000011010, 
18'b000000000000001110, 
18'b111111111111101110, 
18'b111111111110011000, 
18'b111111111110001110, 
18'b000000000010000111, 
18'b111111111101110010, 
18'b000000000000001010, 
18'b111111111111111010, 
18'b000000000000000100, 
18'b000000000000101101, 
18'b111111111111100101, 
18'b000000000000010001, 
18'b111111111111001000, 
18'b000000000000110100, 
18'b111111111111111111, 
18'b000000000001001000, 
18'b000000000000101110, 
18'b111111111111001000, 
18'b000000000000111011, 
18'b000000000000111011, 
18'b000000000000000010, 
18'b000000000000101101, 
18'b111111111111001111, 
18'b111111111101100100, 
18'b111111111111110110, 
18'b111111111110101000, 
18'b111111111111011101, 
18'b000000000000010011, 
18'b000000000001100110, 
18'b000000000000011000, 
18'b000000000000101111, 
18'b111111111111011100, 
18'b000000000000010100, 
18'b000000000000101010, 
18'b111111111111011110, 
18'b000000000000110011, 
18'b000000000001100111, 
18'b000000000000111111, 
18'b000000000000100110, 
18'b111111111111101100, 
18'b000000000000011000, 
18'b000000000001001011, 
18'b000000000000101010, 
18'b111111111110000110, 
18'b000000000000001001, 
18'b111111111111101010, 
18'b111111111111111101, 
18'b000000000001000010, 
18'b111111111101110110, 
18'b111111111110111001, 
18'b000000000000110110, 
18'b000000000001101110, 
18'b000000000000001001, 
18'b000000000001101111, 
18'b111111111101111100, 
18'b000000000000000100, 
18'b000000000000111101, 
18'b000000000010001110, 
18'b111111111101111000, 
18'b111111111111010100, 
18'b111111111101011101, 
18'b111111111111100000, 
18'b000000000000110011, 
18'b111111111110111111, 
18'b000000000000010110, 
18'b111111111111010011, 
18'b111111111110110100, 
18'b000000000000111100, 
18'b111111111111010100, 
18'b111111111111100111, 
18'b111111111110100000, 
18'b000000000000010011, 
18'b111111111111011100, 
18'b000000000000011110, 
18'b111111111111001011, 
18'b000000000001010001, 
18'b111111111110111001, 
18'b000000000001010001, 
18'b111111111111011010, 
18'b111111111101001101, 
18'b000000000000011001, 
18'b000000000001001101, 
18'b000000000000000101, 
18'b000000000000001101, 
18'b000000000000010000, 
18'b000000000001010010, 
18'b111111111111001110, 
18'b000000000000010111, 
18'b111111111110000011, 
18'b000000000001000000, 
18'b000000000001001000, 
18'b000000000000001001, 
18'b111111111111011110, 
18'b000000000000101001, 
18'b111111111111100001, 
18'b000000000000100010, 
18'b000000000000010001, 
18'b000000000000000000, 
18'b000000000000001100, 
18'b111111111110110011, 
18'b000000000000011000, 
18'b111111111111101001, 
18'b000000000000010011, 
18'b000000000001101010, 
18'b000000000001000101, 
18'b111111111111110100, 
18'b111111111110011010, 
18'b000000000000111001, 
18'b111111111110001010, 
18'b111111111111011111, 
18'b111111111111001111, 
18'b111111111111111101, 
18'b000000000001010111, 
18'b111111111111100101, 
18'b000000000000000001, 
18'b000000000001111100, 
18'b111111111111101000, 
18'b111111111111101000, 
18'b111111111111011110, 
18'b111111111111110110, 
18'b000000000001000010, 
18'b111111111110100100, 
18'b111111111111010011, 
18'b111111111111010101, 
18'b111111111110011101, 
18'b111111111110111100, 
18'b111111111101111010, 
18'b111111111111001011, 
18'b111111111111001110, 
18'b111111111101111111, 
18'b000000000001100011, 
18'b111111111110011111, 
18'b000000000000100011, 
18'b111111111110101011, 
18'b111111111110101100, 
18'b000000000000111101, 
18'b000000000000000001, 
18'b111111111110100101, 
18'b000000000000010111, 
18'b111111111110010111, 
18'b000000000001010010, 
18'b000000000000100100, 
18'b111111111111011010, 
18'b111111111110111101, 
18'b111111111111000001, 
18'b000000000000110011, 
18'b111111111110100000, 
18'b000000000000000101, 
18'b000000000001010010, 
18'b000000000000101100, 
18'b000000000000110110, 
18'b111111111110100110, 
18'b000000000001100111, 
18'b000000000001001110, 
18'b000000000000001100, 
18'b000000000001110100, 
18'b000000000000001110, 
18'b111111111101110011, 
18'b000000000001101100, 
18'b000000000000101001, 
18'b000000000001011001, 
18'b111111111110001110, 
18'b111111111111101001, 
18'b000000000000011100, 
18'b111111111110100111, 
18'b111111111110110010, 
18'b111111111110110111, 
18'b111111111111001011, 
18'b000000000001110101, 
18'b000000000000000110, 
18'b000000000000110100, 
18'b000000000000000110, 
18'b000000000001100001, 
18'b000000000001011100, 
18'b111111111110000111, 
18'b111111111110101100, 
18'b000000000001000110, 
18'b111111111110111101, 
18'b111111111111101100, 
18'b111111111111101100, 
18'b000000000001000001, 
18'b000000000000011000, 
18'b111111111111111011, 
18'b111111111110101010, 
18'b000000000001001111, 
18'b111111111111100101, 
18'b000000000001010111, 
18'b000000000000011110, 
18'b000000000000101010, 
18'b111111111111011111, 
18'b000000000000001000, 
18'b000000000001010111, 
18'b111111111111101110, 
18'b111111111111111010, 
18'b111111111111110100, 
18'b111111111110110011, 
18'b000000000010000000, 
18'b000000000000010011, 
18'b111111111111000010, 
18'b111111111111110101, 
18'b000000000000011100, 
18'b111111111111101001, 
18'b111111111111101000, 
18'b000000000000010010, 
18'b000000000001100101, 
18'b000000000000111000, 
18'b000000000001011011, 
18'b000000000000011111, 
18'b111111111110110100, 
18'b000000000000010100, 
18'b111111111110110100, 
18'b111111111111010101, 
18'b111111111111000010, 
18'b000000000000000000, 
18'b000000000000001011, 
18'b000000000000101011, 
18'b000000000000011001, 
18'b000000000000100000, 
18'b111111111101100111, 
18'b111111111110110000, 
18'b111111111111110000, 
18'b000000000000001110, 
18'b000000000001111011, 
18'b000000000001111000, 
18'b111111111101111001, 
18'b111111111111101111, 
18'b000000000001000010, 
18'b000000000001101011, 
18'b111111111101111001, 
18'b111111111110110100, 
18'b000000000000001110, 
18'b000000000001001011, 
18'b111111111111010001, 
18'b111111111111011101, 
18'b111111111111100100, 
18'b111111111111111010, 
18'b000000000001101011, 
18'b000000000001010100, 
18'b111111111111110110, 
18'b111111111111011011, 
18'b000000000001001011, 
18'b000000000000100100, 
18'b000000000001000101, 
18'b111111111111110011, 
18'b111111111111000011, 
18'b111111111111100011, 
18'b111111111111110010, 
18'b111111111110010100, 
18'b000000000000010110, 
18'b111111111110011000, 
18'b000000000000110011, 
18'b111111111111110000, 
18'b111111111111110010, 
18'b000000000001000001, 
18'b000000000000001001, 
18'b111111111111110101, 
18'b000000000000101011, 
18'b000000000000100001, 
18'b000000000000011011, 
18'b000000000000001101, 
18'b000000000000110000, 
18'b111111111110111110, 
18'b000000000010000001, 
18'b000000000000111111, 
18'b111111111101110100, 
18'b000000000000001001, 
18'b111111111110010000, 
18'b111111111110001100, 
18'b111111111101101011, 
18'b111111111111100101, 
18'b111111111111010101, 
18'b111111111111000001, 
18'b000000000000101101, 
18'b000000000000001000, 
18'b111111111110011111, 
18'b000000000000010100, 
18'b111111111111000011, 
18'b111111111111001000, 
18'b111111111111010000, 
18'b111111111111011110, 
18'b111111111111001100, 
18'b000000000000001000, 
18'b111111111111100100, 
18'b000000000001001011, 
18'b111111111111000000, 
18'b000000000000011011, 
18'b000000000000001100, 
18'b000000000000101100, 
18'b000000000001101100, 
18'b000000000000000000, 
18'b111111111110111010, 
18'b111111111111010000, 
18'b000000000000111001, 
18'b000000000001000111, 
18'b111111111101011110, 
18'b000000000000100110, 
18'b000000000000001001, 
18'b111111111101110101, 
18'b000000000001011010, 
18'b111111111111011000, 
18'b000000000000000010, 
18'b111111111110110111, 
18'b000000000001011000, 
18'b000000000000111110, 
18'b111111111101001101, 
18'b000000000001000111, 
18'b000000000000101111, 
18'b000000000000101100, 
18'b000000000010010100, 
18'b000000000000101001, 
18'b000000000001010001, 
18'b111111111110110001, 
18'b000000000000010010, 
18'b111111111111100010, 
18'b000000000000100010, 
18'b000000000001110110, 
18'b000000000000111011, 
18'b111111111101011101, 
18'b000000000001010011, 
18'b111111111111011011, 
18'b000000000000010110, 
18'b111111111110111110, 
18'b111111111110100100, 
18'b000000000000010001, 
18'b000000000000111100, 
18'b000000000000011110, 
18'b111111111111100011, 
18'b111111111101101100, 
18'b000000000000100101, 
18'b000000000000001101, 
18'b000000000001001010, 
18'b000000000000000011, 
18'b000000000000010001, 
18'b000000000001001110, 
18'b000000000001000100, 
18'b111111111111011011, 
18'b000000000000110111, 
18'b111111111110111110, 
18'b111111111110111111, 
18'b111111111111010100, 
18'b000000000001011001, 
18'b111111111111000011, 
18'b111111111110100111, 
18'b000000000000001110, 
18'b000000000000110111, 
18'b000000000001000100, 
18'b111111111111001110, 
18'b111111111101110111, 
18'b111111111101110011, 
18'b000000000000111101, 
18'b000000000000000111, 
18'b000000000001010111, 
18'b000000000001000110, 
18'b000000000000111011, 
18'b000000000001011100, 
18'b111111111111010011, 
18'b111111111111111000, 
18'b000000000000010110, 
18'b000000000000100101, 
18'b000000000001001110, 
18'b000000000001010111, 
18'b000000000001101000, 
18'b111111111110111100, 
18'b000000000000000000, 
18'b000000000001101010, 
18'b000000000001001101, 
18'b000000000001001000, 
18'b111111111111111001, 
18'b111111111110101111, 
18'b111111111111101010, 
18'b111111111111101101, 
18'b111111111110111100, 
18'b111111111110000010, 
18'b000000000001000011, 
18'b000000000000111100, 
18'b000000000001010000, 
18'b000000000000000001, 
18'b111111111111001111, 
18'b111111111111101011, 
18'b111111111111000011, 
18'b000000000000001111, 
18'b000000000000000001, 
18'b000000000001011110, 
18'b000000000000101001, 
18'b111111111101110001, 
18'b111111111110110111, 
18'b111111111110100101, 
18'b111111111111111100, 
18'b111111111110001100, 
18'b111111111111100111, 
18'b111111111111011010, 
18'b000000000000011011, 
18'b000000000000000100, 
18'b000000000000010001, 
18'b111111111101100110, 
18'b111111111111111010, 
18'b000000000001000101, 
18'b000000000001101100, 
18'b111111111111110101, 
18'b111111111110000111, 
18'b000000000000111100, 
18'b111111111111100011, 
18'b000000000001011010, 
18'b111111111111111101, 
18'b111111111101101111, 
18'b111111111111010000, 
18'b000000000000001011, 
18'b111111111110001001, 
18'b111111111111110101, 
18'b000000000001011010, 
18'b111111111111011010, 
18'b111111111111111010, 
18'b000000000001010111, 
18'b000000000000011101, 
18'b111111111111011011, 
18'b000000000001011100, 
18'b111111111111011100, 
18'b000000000000100110, 
18'b000000000000000110, 
18'b111111111110011101, 
18'b000000000001010000, 
18'b111111111111001101, 
18'b000000000000000100, 
18'b000000000000001010, 
18'b111111111111010011, 
18'b111111111111100110, 
18'b000000000000111000, 
18'b000000000000000001, 
18'b000000000000010110, 
18'b000000000000100110, 
18'b111111111111000111, 
18'b000000000000011101, 
18'b111111111110101011, 
18'b111111111111111101, 
18'b111111111111001101, 
18'b111111111111001010, 
18'b111111111110110010, 
18'b000000000000001100, 
18'b000000000000101010, 
18'b000000000000010111, 
18'b111111111111011000, 
18'b111111111110110101, 
18'b000000000001010100, 
18'b111111111111001111, 
18'b000000000000000000, 
18'b000000000001100111, 
18'b000000000000000010, 
18'b111111111110011001, 
18'b000000000001000110, 
18'b111111111110111001, 
18'b000000000000101110, 
18'b000000000000011111, 
18'b000000000000100000, 
18'b000000000001000011, 
18'b111111111110110000, 
18'b000000000000011001, 
18'b111111111111001100, 
18'b111111111110100010, 
18'b000000000000110111, 
18'b111111111110011101, 
18'b000000000001011010, 
18'b000000000000010001, 
18'b111111111111011100, 
18'b111111111110011001, 
18'b111111111111010011, 
18'b000000000001010100, 
18'b111111111111000001, 
18'b000000000000000101, 
18'b111111111111010100, 
18'b000000000001100000, 
18'b111111111111101111, 
18'b000000000000001001, 
18'b000000000000110000, 
18'b111111111111001101, 
18'b111111111111000110, 
18'b000000000000011000, 
18'b000000000000001100, 
18'b111111111110001010, 
18'b000000000001101101, 
18'b111111111111101001, 
18'b000000000001100101, 
18'b000000000000111000, 
18'b000000000000110010, 
18'b111111111110111000, 
18'b111111111111101000, 
18'b111111111111101000, 
18'b111111111111011100, 
18'b111111111111110101, 
18'b000000000000111000, 
18'b111111111111000001, 
18'b000000000000110011, 
18'b000000000000001011, 
18'b000000000000010001, 
18'b000000000000110100, 
18'b000000000001010000, 
18'b000000000000101010, 
18'b111111111111000100, 
18'b000000000000011101, 
18'b111111111110000111, 
18'b000000000000100010, 
18'b111111111111011010, 
18'b000000000000110001, 
18'b111111111111010010, 
18'b111111111111001001, 
18'b000000000000101010, 
18'b111111111110110001, 
18'b111111111111001111, 
18'b111111111110101001, 
18'b000000000000001110, 
18'b111111111111000110, 
18'b000000000001110011, 
18'b111111111111110100, 
18'b111111111111000100, 
18'b111111111111111110, 
18'b000000000000101001, 
18'b000000000000101000, 
18'b000000000001010111, 
18'b111111111111010111, 
18'b111111111110100000, 
18'b000000000000000110, 
18'b111111111110111101, 
18'b111111111111010111, 
18'b111111111110010000, 
18'b000000000000110110, 
18'b000000000010000110, 
18'b000000000000110011, 
18'b000000000001010011, 
18'b111111111111111100, 
18'b111111111111000110, 
18'b000000000001001000, 
18'b111111111111100001, 
18'b000000000001010001, 
18'b111111111111011001, 
18'b000000000000010111, 
18'b111111111110100011, 
18'b000000000010001100, 
18'b000000000001111001, 
18'b111111111111001001, 
18'b111111111101011100, 
18'b000000000000001011, 
18'b111111111110110001, 
18'b000000000010000001, 
18'b111111111111110000, 
18'b111111111111001101, 
18'b000000000000001101, 
18'b111111111111000110, 
18'b111111111111001010, 
18'b111111111111011101, 
18'b111111111101100111, 
18'b000000000000001111, 
18'b111111111101101010, 
18'b111111111111010101, 
18'b000000000000001101, 
18'b000000000000101110, 
18'b111111111111000111, 
18'b111111111111110111, 
18'b000000000000010100, 
18'b111111111111011011, 
18'b111111111101010100, 
18'b111111111111011010, 
18'b000000000000011010, 
18'b000000000000010010, 
18'b000000000000100101, 
18'b000000000000101000, 
18'b111111111101110111, 
18'b111111111111010000, 
18'b000000000001011000, 
18'b111111111110011100, 
18'b111111111111011100, 
18'b000000000001110111, 
18'b111111111111001100, 
18'b000000000000000011, 
18'b111111111111001110, 
18'b000000000000010000, 
18'b111111111111101011, 
18'b111111111111011100, 
18'b000000000001011111, 
18'b111111111110011111, 
18'b111111111111011100, 
18'b000000000001001001, 
18'b000000000001011101, 
18'b111111111111100101, 
18'b000000000000100001, 
18'b111111111111101100, 
18'b111111111101110100, 
18'b111111111111011110, 
18'b000000000000010010, 
18'b111111111111001110, 
18'b111111111111111100, 
18'b111111111111100000, 
18'b111111111111001110, 
18'b000000000001001101, 
18'b111111111111001110, 
18'b111111111111000000, 
18'b000000000000000110, 
18'b111111111111100000, 
18'b000000000000101000, 
18'b111111111110101100, 
18'b000000000001010000, 
18'b000000000000111111, 
18'b000000000000000101, 
18'b111111111111111101, 
18'b111111111110111000, 
18'b111111111110101011, 
18'b111111111111000110, 
18'b111111111111011011, 
18'b111111111111101111, 
18'b000000000000010100, 
18'b000000000001111001, 
18'b111111111111011101, 
18'b111111111110001110, 
18'b000000000001110101, 
18'b111111111111000110, 
18'b111111111111110010, 
18'b000000000000010001, 
18'b000000000000110101, 
18'b111111111110111110, 
18'b111111111111000100, 
18'b111111111111100110, 
18'b000000000000111011, 
18'b111111111111001110, 
18'b000000000000110010, 
18'b000000000000111010, 
18'b111111111110100110, 
18'b000000000000000011, 
18'b000000000000000001, 
18'b111111111111100110, 
18'b111111111111011001, 
18'b000000000000001011, 
18'b111111111111100111, 
18'b000000000000011100, 
18'b000000000000011011, 
18'b111111111110101001, 
18'b111111111111000100, 
18'b000000000000001110, 
18'b000000000000111100, 
18'b111111111110010000, 
18'b111111111101110011, 
18'b111111111111001110, 
18'b111111111111101001, 
18'b111111111111101111, 
18'b111111111111110110, 
18'b111111111110110110, 
18'b000000000000101011, 
18'b000000000000101111, 
18'b111111111111001110, 
18'b000000000000110110, 
18'b111111111111111000, 
18'b111111111111011101, 
18'b000000000001011000, 
18'b111111111111000011, 
18'b111111111111101101, 
18'b111111111111000011, 
18'b000000000000011001, 
18'b000000000001001000, 
18'b111111111111111100, 
18'b000000000000101101, 
18'b111111111101101110, 
18'b000000000000001101, 
18'b111111111111001011, 
18'b111111111111010110, 
18'b000000000001001101, 
18'b111111111110100011, 
18'b000000000000101010, 
18'b111111111111010111, 
18'b000000000000000010, 
18'b000000000000000010, 
18'b111111111110011001, 
18'b111111111111111001, 
18'b000000000000001111, 
18'b111111111110110110, 
18'b000000000000010000, 
18'b000000000001010000, 
18'b111111111111001000, 
18'b000000000000111100, 
18'b111111111111100011, 
18'b000000000001101111, 
18'b111111111101011111, 
18'b111111111101011000, 
18'b000000000000110001, 
18'b111111111111010010, 
18'b000000000000010101, 
18'b111111111110111011, 
18'b111111111111101011, 
18'b000000000000111011, 
18'b000000000000010001, 
18'b111111111111111100, 
18'b000000000000010000, 
18'b111111111111001001, 
18'b000000000001000101, 
18'b111111111111111101, 
18'b111111111111001110, 
18'b000000000000101000, 
18'b111111111111110001, 
18'b000000000000000111, 
18'b000000000000111110, 
18'b111111111110010011, 
18'b111111111111000000, 
18'b111111111101011110, 
18'b000000000000100000, 
18'b111111111110010010, 
18'b000000000000110000, 
18'b000000000000100111, 
18'b111111111111111111, 
18'b111111111110111111, 
18'b111111111111001011, 
18'b000000000000111001, 
18'b111111111111110100, 
18'b111111111101111110, 
18'b000000000001100101, 
18'b111111111101110001, 
18'b111111111110110011, 
18'b111111111111110000, 
18'b000000000000000000, 
18'b111111111110100100, 
18'b111111111111010110, 
18'b111111111111111110, 
18'b111111111111110110, 
18'b111111111111101000, 
18'b111111111111111010, 
18'b111111111111000101, 
18'b000000000001110001, 
18'b111111111111100010, 
18'b000000000000001110, 
18'b000000000000001110, 
18'b111111111111101100, 
18'b000000000000010100, 
18'b000000000000001011, 
18'b111111111111100111, 
18'b111111111111101001, 
18'b000000000000011011, 
18'b000000000000001101, 
18'b000000000000010110, 
18'b000000000000101011, 
18'b111111111110110100, 
18'b000000000001111100, 
18'b111111111111010000, 
18'b000000000000010000, 
18'b111111111111010100, 
18'b000000000000101001, 
18'b111111111110100111, 
18'b111111111110111001, 
18'b111111111110001110, 
18'b111111111111101010, 
18'b111111111101011001, 
18'b111111111111111011, 
18'b111111111111000111, 
18'b111111111110100100, 
18'b111111111110111100, 
18'b111111111111011111, 
18'b111111111111000100, 
18'b000000000001010100, 
18'b111111111101011110, 
18'b000000000010000100, 
18'b111111111111101011, 
18'b111111111110111101, 
18'b111111111111101010, 
18'b111111111110011101, 
18'b000000000000010010, 
18'b000000000000101100, 
18'b111111111110101011, 
18'b000000000000010111, 
18'b111111111110001001, 
18'b000000000001000010, 
18'b111111111110011111, 
18'b000000000000010111, 
18'b111111111111010001, 
18'b111111111111100001, 
18'b000000000001011001, 
18'b000000000001001001, 
18'b111111111111001100, 
18'b000000000001000111, 
18'b000000000000011100, 
18'b000000000000010011, 
18'b000000000001101101, 
18'b000000000000111110, 
18'b111111111111001000, 
18'b111111111111000000, 
18'b000000000001011100, 
18'b000000000001010101, 
18'b000000000000000111, 
18'b000000000000110000, 
18'b000000000000010111, 
18'b000000000000010110, 
18'b111111111111101100, 
18'b000000000001001111, 
18'b111111111111110000, 
18'b000000000000000001, 
18'b000000000000011110, 
18'b000000000010011001, 
18'b111111111110101011, 
18'b111111111111011101, 
18'b000000000000000011, 
18'b000000000001000000, 
18'b000000000001001111, 
18'b111111111110110001, 
18'b111111111110101100, 
18'b000000000000001010, 
18'b000000000000011100, 
18'b000000000000001010, 
18'b000000000000010000, 
18'b000000000000100100, 
18'b000000000000011101, 
18'b000000000001000010, 
18'b111111111111111100, 
18'b000000000000001011, 
18'b000000000001001000, 
18'b111111111111111011, 
18'b111111111111101000, 
18'b000000000000010000, 
18'b111111111110011001, 
18'b000000000000001100, 
18'b000000000000101100, 
18'b111111111110101110, 
18'b000000000001111101, 
18'b111111111111111000, 
18'b000000000000011111, 
18'b111111111111111010, 
18'b111111111111101101, 
18'b111111111111101001, 
18'b000000000000111011, 
18'b000000000001111110, 
18'b000000000000000000, 
18'b000000000000110000, 
18'b000000000010000001, 
18'b111111111110011110, 
18'b000000000000111100, 
18'b000000000001000001, 
18'b111111111110111101, 
18'b000000000000001111, 
18'b000000000001001110, 
18'b000000000000000111, 
18'b000000000000111010, 
18'b111111111111110111, 
18'b000000000001101110, 
18'b000000000000101111, 
18'b111111111111010001, 
18'b111111111110000111, 
18'b111111111110110111, 
18'b000000000000011001, 
18'b000000000000000111, 
18'b111111111111110000, 
18'b000000000000100011, 
18'b000000000000101101, 
18'b000000000000101010, 
18'b111111111110001100, 
18'b000000000000010111, 
18'b000000000000110100, 
18'b111111111110011011, 
18'b111111111111001011, 
18'b111111111111101110, 
18'b000000000001100100, 
18'b000000000001101010, 
18'b111111111111111110, 
18'b000000000000111010, 
18'b111111111110011010, 
18'b111111111111011010, 
18'b111111111111011110, 
18'b111111111111110010, 
18'b000000000000001001, 
18'b111111111101111000, 
18'b000000000000111011, 
18'b111111111111100101, 
18'b111111111111100100, 
18'b111111111110101000, 
18'b000000000000001110, 
18'b111111111111111011, 
18'b000000000010010111, 
18'b111111111110001011, 
18'b000000000000100000, 
18'b000000000000000011, 
18'b111111111111000010, 
18'b111111111111011001, 
18'b000000000000010100, 
18'b111111111110101011, 
18'b111111111111001110, 
18'b111111111110001111, 
18'b111111111111100011, 
18'b000000000000110111, 
18'b000000000001100110, 
18'b111111111110111101, 
18'b111111111111100110, 
18'b000000000000010011, 
18'b000000000001010010, 
18'b111111111111011110, 
18'b111111111111111110, 
18'b111111111111110101, 
18'b000000000001011000, 
18'b111111111101110111, 
18'b000000000001010101, 
18'b111111111111001000, 
18'b111111111101111100, 
18'b111111111110111100, 
18'b000000000010000101, 
18'b111111111110010111, 
18'b111111111111100010, 
18'b111111111110000001, 
18'b000000000000110001, 
18'b000000000001110000, 
18'b000000000001110110, 
18'b111111111110111110, 
18'b000000000000000110, 
18'b111111111101111001, 
18'b000000000000110110, 
18'b111111111111000010, 
18'b000000000001001011, 
18'b000000000000000010, 
18'b000000000000101000, 
18'b111111111111000001, 
18'b111111111111001101, 
18'b111111111110111011, 
18'b000000000000011001, 
18'b000000000000100011, 
18'b000000000001101111, 
18'b000000000000010001, 
18'b111111111111000010, 
18'b111111111111100001, 
18'b111111111110010010, 
18'b000000000001010101, 
18'b000000000000111011, 
18'b111111111110100010, 
18'b111111111111100111, 
18'b111111111101111001, 
18'b000000000001010101, 
18'b111111111110011001, 
18'b000000000001101000, 
18'b111111111110111111, 
18'b000000000000011000, 
18'b000000000000001101, 
18'b000000000001010000, 
18'b111111111110110111, 
18'b111111111110101111, 
18'b000000000001011010, 
18'b111111111111001101, 
18'b000000000000001010, 
18'b111111111110101010, 
18'b000000000000000110, 
18'b111111111111010000, 
18'b000000000000111010, 
18'b111111111111011010, 
18'b111111111111001101, 
18'b111111111111010000, 
18'b000000000000110010, 
18'b111111111111011001, 
18'b111111111111101010, 
18'b000000000000101000, 
18'b000000000001001101, 
18'b111111111110000101, 
18'b000000000000001001, 
18'b000000000000001101, 
18'b111111111101111100, 
18'b111111111111101100, 
18'b000000000001100010, 
18'b000000000000111010, 
18'b111111111110001110, 
18'b000000000000111101, 
18'b111111111100100010, 
18'b111111111110010111, 
18'b111111111110100101, 
18'b000000000000001000, 
18'b111111111101110101, 
18'b111111111111011100, 
18'b000000000000001001, 
18'b111111111111010000, 
18'b000000000001111111, 
18'b000000000000010000, 
18'b000000000000000101, 
18'b000000000000000000, 
18'b000000000010010110, 
18'b111111111110100111, 
18'b111111111110101111, 
18'b000000000000010111, 
18'b000000000001010100, 
18'b000000000001000000, 
18'b000000000001000001, 
18'b111111111111000101, 
18'b111111111110101111, 
18'b000000000000001111, 
18'b111111111110111010, 
18'b000000000000010101, 
18'b000000000000011111, 
18'b000000000000001010, 
18'b111111111110001011, 
18'b111111111110001010, 
18'b111111111111110010, 
18'b111111111111100011, 
18'b111111111111101101, 
18'b111111111110000010, 
18'b000000000000010101, 
18'b111111111111010100, 
18'b111111111101101010, 
18'b111111111110111101, 
18'b000000000001010111, 
18'b111111111110011110, 
18'b000000000001001001, 
18'b000000000010000001, 
18'b000000000001111110, 
18'b111111111111111100, 
18'b111111111110101011, 
18'b000000000000110111, 
18'b111111111110101100, 
18'b111111111111011100, 
18'b000000000000110011, 
18'b111111111111110010, 
18'b111111111111101111, 
18'b111111111111101101, 
18'b000000000001000001 

};
localparam logic signed [17:0] dlBiases [9:0] = {
18'b000000000001010101, 
18'b111111111111111111, 
18'b111111111111111111, 
18'b111111111111100010, 
18'b111111111111100000, 
18'b111111111111110101, 
18'b111111111111110100, 
18'b000000000000100111, 
18'b111111111110100011, 
18'b111111111111110101

};
localparam logic signed [17:0] convWeights [0:17] = {
18'b000000000000111001, 
18'b000000000011110110, 
18'b111111111110000101, 
18'b000000000000101111, 
18'b000000000000000111, 
18'b000000000100000110, 
18'b000000000011001111, 
18'b000000000001100110, 
18'b111111111110001011, 
18'b000000000010110010, 
18'b111111111111010011, 
18'b000000000001101011, 
18'b000000000011111110, 
18'b000000000001010001, 
18'b000000000011000100, 
18'b111111111111111010, 
18'b000000000001011101, 
18'b000000000000111010

};
localparam logic signed [17:0] convBiases [1:0] = {
18'b000000000000000000, 
18'b000000000000000000

};
endpackage